
module decode
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  input_r,
  ih_i,
  ih_o,
  ih_o_ap_vld,
  dec_del_bpl_address0,
  dec_del_bpl_ce0,
  dec_del_bpl_we0,
  dec_del_bpl_d0,
  dec_del_bpl_q0,
  dec_del_dltx_address0,
  dec_del_dltx_ce0,
  dec_del_dltx_we0,
  dec_del_dltx_d0,
  dec_del_dltx_q0,
  dec_del_dltx_address1,
  dec_del_dltx_ce1,
  dec_del_dltx_we1,
  dec_del_dltx_d1,
  dec_del_dltx_q1,
  dec_rlt1_i,
  dec_rlt1_o,
  dec_rlt1_o_ap_vld,
  dec_al1_i,
  dec_al1_o,
  dec_al1_o_ap_vld,
  dec_rlt2_i,
  dec_rlt2_o,
  dec_rlt2_o_ap_vld,
  dec_al2_i,
  dec_al2_o,
  dec_al2_o_ap_vld,
  dec_detl_i,
  dec_detl_o,
  dec_detl_o_ap_vld,
  il,
  dec_nbl_i,
  dec_nbl_o,
  dec_nbl_o_ap_vld,
  dec_plt1_i,
  dec_plt1_o,
  dec_plt1_o_ap_vld,
  dec_plt2_i,
  dec_plt2_o,
  dec_plt2_o_ap_vld,
  dec_del_bph_address0,
  dec_del_bph_ce0,
  dec_del_bph_we0,
  dec_del_bph_d0,
  dec_del_bph_q0,
  dec_del_dhx_address0,
  dec_del_dhx_ce0,
  dec_del_dhx_we0,
  dec_del_dhx_d0,
  dec_del_dhx_q0,
  dec_del_dhx_address1,
  dec_del_dhx_ce1,
  dec_del_dhx_we1,
  dec_del_dhx_d1,
  dec_del_dhx_q1,
  dec_rh1_i,
  dec_rh1_o,
  dec_rh1_o_ap_vld,
  dec_ah1_i,
  dec_ah1_o,
  dec_ah1_o_ap_vld,
  dec_rh2_i,
  dec_rh2_o,
  dec_rh2_o_ap_vld,
  dec_ah2_i,
  dec_ah2_o,
  dec_ah2_o_ap_vld,
  dec_deth_i,
  dec_deth_o,
  dec_deth_o_ap_vld,
  dec_nbh_i,
  dec_nbh_o,
  dec_nbh_o_ap_vld,
  dec_ph1_i,
  dec_ph1_o,
  dec_ph1_o_ap_vld,
  dec_ph2_i,
  dec_ph2_o,
  dec_ph2_o_ap_vld,
  accumc_address0,
  accumc_ce0,
  accumc_we0,
  accumc_d0,
  accumc_q0,
  accumd_address0,
  accumd_ce0,
  accumd_we0,
  accumd_d0,
  accumd_q0,
  working_key
);

  parameter ap_ST_fsm_state1 = 29'd1;
  parameter ap_ST_fsm_state2 = 29'd2;
  parameter ap_ST_fsm_state3 = 29'd4;
  parameter ap_ST_fsm_state4 = 29'd8;
  parameter ap_ST_fsm_state5 = 29'd16;
  parameter ap_ST_fsm_state6 = 29'd32;
  parameter ap_ST_fsm_state7 = 29'd64;
  parameter ap_ST_fsm_state8 = 29'd128;
  parameter ap_ST_fsm_state9 = 29'd256;
  parameter ap_ST_fsm_state10 = 29'd512;
  parameter ap_ST_fsm_state11 = 29'd1024;
  parameter ap_ST_fsm_state12 = 29'd2048;
  parameter ap_ST_fsm_state13 = 29'd4096;
  parameter ap_ST_fsm_state14 = 29'd8192;
  parameter ap_ST_fsm_state15 = 29'd16384;
  parameter ap_ST_fsm_state16 = 29'd32768;
  parameter ap_ST_fsm_state17 = 29'd65536;
  parameter ap_ST_fsm_state18 = 29'd131072;
  parameter ap_ST_fsm_state19 = 29'd262144;
  parameter ap_ST_fsm_state20 = 29'd524288;
  parameter ap_ST_fsm_state21 = 29'd1048576;
  parameter ap_ST_fsm_state22 = 29'd2097152;
  parameter ap_ST_fsm_state23 = 29'd4194304;
  parameter ap_ST_fsm_state24 = 29'd8388608;
  parameter ap_ST_fsm_state25 = 29'd16777216;
  parameter ap_ST_fsm_state26 = 29'd33554432;
  parameter ap_ST_fsm_state27 = 29'd67108864;
  parameter ap_ST_fsm_state28 = 29'd134217728;
  parameter ap_ST_fsm_state29 = 29'd268435456;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  input [31:0] input_r;
  input [31:0] ih_i;
  output [31:0] ih_o;
  output ih_o_ap_vld;
  output [2:0] dec_del_bpl_address0;
  output dec_del_bpl_ce0;
  output dec_del_bpl_we0;
  output [31:0] dec_del_bpl_d0;
  input [31:0] dec_del_bpl_q0;
  output [2:0] dec_del_dltx_address0;
  output dec_del_dltx_ce0;
  output dec_del_dltx_we0;
  output [31:0] dec_del_dltx_d0;
  input [31:0] dec_del_dltx_q0;
  output [2:0] dec_del_dltx_address1;
  output dec_del_dltx_ce1;
  output dec_del_dltx_we1;
  output [31:0] dec_del_dltx_d1;
  input [31:0] dec_del_dltx_q1;
  input [31:0] dec_rlt1_i;
  output [31:0] dec_rlt1_o;
  output dec_rlt1_o_ap_vld;
  input [31:0] dec_al1_i;
  output [31:0] dec_al1_o;
  output dec_al1_o_ap_vld;
  input [31:0] dec_rlt2_i;
  output [31:0] dec_rlt2_o;
  output dec_rlt2_o_ap_vld;
  input [31:0] dec_al2_i;
  output [31:0] dec_al2_o;
  output dec_al2_o_ap_vld;
  input [14:0] dec_detl_i;
  output [14:0] dec_detl_o;
  output dec_detl_o_ap_vld;
  input [5:0] il;
  input [31:0] dec_nbl_i;
  output [31:0] dec_nbl_o;
  output dec_nbl_o_ap_vld;
  input [31:0] dec_plt1_i;
  output [31:0] dec_plt1_o;
  output dec_plt1_o_ap_vld;
  input [31:0] dec_plt2_i;
  output [31:0] dec_plt2_o;
  output dec_plt2_o_ap_vld;
  output [2:0] dec_del_bph_address0;
  output dec_del_bph_ce0;
  output dec_del_bph_we0;
  output [31:0] dec_del_bph_d0;
  input [31:0] dec_del_bph_q0;
  output [2:0] dec_del_dhx_address0;
  output dec_del_dhx_ce0;
  output dec_del_dhx_we0;
  output [31:0] dec_del_dhx_d0;
  input [31:0] dec_del_dhx_q0;
  output [2:0] dec_del_dhx_address1;
  output dec_del_dhx_ce1;
  output dec_del_dhx_we1;
  output [31:0] dec_del_dhx_d1;
  input [31:0] dec_del_dhx_q1;
  input [31:0] dec_rh1_i;
  output [31:0] dec_rh1_o;
  output dec_rh1_o_ap_vld;
  input [31:0] dec_ah1_i;
  output [31:0] dec_ah1_o;
  output dec_ah1_o_ap_vld;
  input [31:0] dec_rh2_i;
  output [31:0] dec_rh2_o;
  output dec_rh2_o_ap_vld;
  input [31:0] dec_ah2_i;
  output [31:0] dec_ah2_o;
  output dec_ah2_o_ap_vld;
  input [14:0] dec_deth_i;
  output [14:0] dec_deth_o;
  output dec_deth_o_ap_vld;
  input [31:0] dec_nbh_i;
  output [31:0] dec_nbh_o;
  output dec_nbh_o_ap_vld;
  input [31:0] dec_ph1_i;
  output [31:0] dec_ph1_o;
  output dec_ph1_o_ap_vld;
  input [31:0] dec_ph2_i;
  output [31:0] dec_ph2_o;
  output dec_ph2_o_ap_vld;
  output [3:0] accumc_address0;
  output accumc_ce0;
  output accumc_we0;
  output [31:0] accumc_d0;
  input [31:0] accumc_q0;
  output [3:0] accumd_address0;
  output accumd_ce0;
  output accumd_we0;
  output [31:0] accumd_d0;
  input [31:0] accumd_q0;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [31:0] ih_o;
  reg ih_o_ap_vld;
  reg [2:0] dec_del_bpl_address0;
  reg dec_del_bpl_ce0;
  reg dec_del_bpl_we0;
  reg [2:0] dec_del_dltx_address0;
  reg dec_del_dltx_ce0;
  reg dec_del_dltx_we0;
  reg dec_del_dltx_ce1;
  reg dec_del_dltx_we1;
  reg [31:0] dec_rlt1_o;
  reg dec_rlt1_o_ap_vld;
  reg [31:0] dec_al1_o;
  reg dec_al1_o_ap_vld;
  reg [31:0] dec_rlt2_o;
  reg dec_rlt2_o_ap_vld;
  reg [31:0] dec_al2_o;
  reg dec_al2_o_ap_vld;
  reg [14:0] dec_detl_o;
  reg dec_detl_o_ap_vld;
  reg [31:0] dec_nbl_o;
  reg dec_nbl_o_ap_vld;
  reg [31:0] dec_plt1_o;
  reg dec_plt1_o_ap_vld;
  reg [31:0] dec_plt2_o;
  reg dec_plt2_o_ap_vld;
  reg [2:0] dec_del_bph_address0;
  reg dec_del_bph_ce0;
  reg dec_del_bph_we0;
  reg [2:0] dec_del_dhx_address0;
  reg dec_del_dhx_ce0;
  reg dec_del_dhx_we0;
  reg dec_del_dhx_ce1;
  reg dec_del_dhx_we1;
  reg [31:0] dec_rh1_o;
  reg dec_rh1_o_ap_vld;
  reg [31:0] dec_ah1_o;
  reg dec_ah1_o_ap_vld;
  reg [31:0] dec_rh2_o;
  reg dec_rh2_o_ap_vld;
  reg [31:0] dec_ah2_o;
  reg dec_ah2_o_ap_vld;
  reg [14:0] dec_deth_o;
  reg dec_deth_o_ap_vld;
  reg [31:0] dec_nbh_o;
  reg dec_nbh_o_ap_vld;
  reg [31:0] dec_ph1_o;
  reg dec_ph1_o_ap_vld;
  reg [31:0] dec_ph2_o;
  reg dec_ph2_o_ap_vld;
  reg [3:0] accumc_address0;
  reg accumc_ce0;
  reg accumc_we0;
  reg [31:0] accumc_d0;
  reg [3:0] accumd_address0;
  reg accumd_ce0;
  reg accumd_we0;
  reg [31:0] accumd_d0;
  reg [28:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  wire [3:0] qq4_code4_table_address0;
  reg qq4_code4_table_ce0;
  wire [15:0] qq4_code4_table_q0;
  reg [31:0] dec_dlt;
  wire [5:0] qq6_code6_table_address0;
  reg qq6_code6_table_ce0;
  wire [15:0] qq6_code6_table_q0;
  wire [3:0] wl_code_table_address0;
  reg wl_code_table_ce0;
  wire [12:0] wl_code_table_q0;
  reg [4:0] ilb_table_address0;
  reg ilb_table_ce0;
  wire [11:0] ilb_table_q0;
  reg [31:0] dec_plt;
  reg [31:0] dec_dh;
  reg [31:0] dec_ph;
  reg signed [31:0] reg_477;
  wire ap_CS_fsm_state2;
  wire ap_CS_fsm_state6;
  reg signed [31:0] reg_481;
  reg signed [31:0] reg_485;
  wire ap_CS_fsm_state14;
  wire ap_CS_fsm_state18;
  reg signed [31:0] reg_489;
  wire [31:0] zl_fu_499_p2;
  reg [31:0] zl_reg_1885;
  wire ap_CS_fsm_state3;
  wire ap_CS_fsm_state4;
  wire [2:0] p_01_rec_i_fu_539_p2;
  reg [2:0] p_01_rec_i_reg_1895;
  wire ap_CS_fsm_state5;
  wire [0:0] exitcond3_fu_551_p2;
  wire [31:0] tmp_i_fu_581_p2;
  reg [31:0] tmp_i_reg_1928;
  wire ap_CS_fsm_state7;
  wire [31:0] zl_5_fu_587_p2;
  wire ap_CS_fsm_state8;
  reg signed [15:0] qq4_code4_table_load_reg_1938;
  wire ap_CS_fsm_state9;
  reg signed [15:0] qq6_code6_table_load_reg_1943;
  wire [24:0] nbl_assign_4_cast_fu_636_p2;
  reg [24:0] nbl_assign_4_cast_reg_1948;
  reg [0:0] tmp_73_reg_1953;
  wire [31:0] pl_fu_654_p2;
  reg [31:0] pl_reg_1958;
  wire ap_CS_fsm_state10;
  wire [31:0] tmp_i1_fu_660_p2;
  reg [31:0] tmp_i1_reg_1963;
  wire signed [15:0] tmp_70_fu_677_p4;
  reg signed [15:0] tmp_70_reg_1968;
  reg [15:0] tmp_71_reg_1974;
  reg [3:0] wd2_cast_reg_1979;
  wire signed [16:0] tmp_43_fu_809_p1;
  reg signed [16:0] tmp_43_reg_1989;
  wire ap_CS_fsm_state11;
  wire [18:0] rl_fu_819_p2;
  reg [18:0] rl_reg_1994;
  wire [31:0] tmp_i8_fu_904_p2;
  reg [31:0] tmp_i8_reg_1999;
  wire ap_CS_fsm_state12;
  wire grp_upzero_fu_442_ap_ready;
  wire grp_upzero_fu_442_ap_done;
  wire [31:0] tmp_5_i_fu_910_p2;
  reg [31:0] tmp_5_i_reg_2004;
  reg [0:0] tmp_81_reg_2009;
  wire [26:0] apl2_fu_1038_p2;
  reg [26:0] apl2_reg_2014;
  wire ap_CS_fsm_state13;
  reg [23:0] tmp_21_i_reg_2020;
  wire signed [14:0] apl2_assign_fu_1088_p3;
  reg signed [14:0] apl2_assign_reg_2025;
  wire [24:0] apl1_fu_1112_p2;
  reg [24:0] apl1_reg_2031;
  wire [15:0] tmp_82_fu_1152_p1;
  reg [15:0] tmp_82_reg_2037;
  wire ap_CS_fsm_state15;
  wire signed [15:0] apl1_11_fu_1156_p2;
  reg signed [15:0] apl1_11_reg_2042;
  wire [0:0] tmp_7_i_fu_1166_p2;
  reg [0:0] tmp_7_i_reg_2047;
  wire [31:0] grp_fu_493_p2;
  reg [31:0] zl_4_reg_2052;
  wire signed [31:0] rl_cast_fu_1172_p1;
  reg signed [31:0] rl_cast_reg_2057;
  wire ap_CS_fsm_state16;
  wire [2:0] p_01_rec_i2_fu_1190_p2;
  reg [2:0] p_01_rec_i2_reg_2063;
  wire ap_CS_fsm_state17;
  wire signed [31:0] tmp_14_fu_1216_p6;
  reg signed [31:0] tmp_14_reg_2081;
  wire [0:0] exitcond2_fu_1202_p2;
  wire [30:0] nbh_assign_2_cast_fu_1288_p2;
  reg [30:0] nbh_assign_2_cast_reg_2086;
  reg [0:0] tmp_86_reg_2091;
  reg [31:0] tmp_i8_33_reg_2096;
  wire ap_CS_fsm_state19;
  wire [31:0] zl_6_fu_1302_p2;
  wire ap_CS_fsm_state20;
  reg signed [16:0] tmp_50_reg_2106;
  wire ap_CS_fsm_state21;
  reg [3:0] wd2_17_cast_reg_2113;
  wire signed [18:0] tmp_i19_cast_fu_1399_p1;
  reg signed [18:0] tmp_i19_cast_reg_2123;
  wire ap_CS_fsm_state22;
  wire [31:0] tmp_i3_fu_1472_p2;
  reg [31:0] tmp_i3_reg_2128;
  wire ap_CS_fsm_state23;
  wire [31:0] tmp_5_i5_fu_1478_p2;
  reg [31:0] tmp_5_i5_reg_2133;
  reg [0:0] tmp_94_reg_2138;
  wire [26:0] apl2_2_fu_1606_p2;
  reg [26:0] apl2_2_reg_2143;
  wire ap_CS_fsm_state24;
  reg [23:0] tmp_21_i2_reg_2149;
  wire [31:0] pl_2_fu_1638_p2;
  reg [31:0] pl_2_reg_2154;
  wire ap_CS_fsm_state25;
  wire [31:0] tmp_i4_fu_1644_p2;
  reg [31:0] tmp_i4_reg_2159;
  wire signed [14:0] apl2_assign_2_fu_1672_p3;
  reg signed [14:0] apl2_assign_2_reg_2164;
  wire [24:0] apl1_13_fu_1696_p2;
  reg [24:0] apl1_13_reg_2170;
  wire [15:0] tmp_95_fu_1754_p1;
  reg [15:0] tmp_95_reg_2176;
  wire ap_CS_fsm_state26;
  wire signed [15:0] apl1_15_fu_1758_p2;
  reg signed [15:0] apl1_15_reg_2181;
  wire [0:0] tmp_7_i2_fu_1768_p2;
  reg [0:0] tmp_7_i2_reg_2186;
  wire [18:0] tmp8_fu_1774_p2;
  reg [18:0] tmp8_reg_2191;
  wire [31:0] xd_fu_1819_p2;
  reg [31:0] xd_reg_2196;
  wire ap_CS_fsm_state27;
  wire [31:0] xs_fu_1824_p2;
  reg [31:0] xs_reg_2201;
  reg [3:0] accumc_addr_reg_2206;
  wire ap_CS_fsm_state28;
  reg [3:0] accumd_addr_reg_2211;
  wire [4:0] p_rec_fu_1841_p2;
  reg [4:0] p_rec_reg_2216;
  wire [3:0] i_fu_1865_p2;
  reg [3:0] i_reg_2234;
  wire grp_upzero_fu_442_ap_start;
  wire grp_upzero_fu_442_ap_idle;
  reg [16:0] grp_upzero_fu_442_dlt;
  wire [2:0] grp_upzero_fu_442_dlti_address0;
  wire grp_upzero_fu_442_dlti_ce0;
  wire grp_upzero_fu_442_dlti_we0;
  wire [31:0] grp_upzero_fu_442_dlti_d0;
  reg [31:0] grp_upzero_fu_442_dlti_q0;
  wire [2:0] grp_upzero_fu_442_dlti_address1;
  wire grp_upzero_fu_442_dlti_ce1;
  wire grp_upzero_fu_442_dlti_we1;
  wire [31:0] grp_upzero_fu_442_dlti_d1;
  reg [31:0] grp_upzero_fu_442_dlti_q1;
  wire [2:0] grp_upzero_fu_442_bli_address0;
  wire grp_upzero_fu_442_bli_ce0;
  wire grp_upzero_fu_442_bli_we0;
  wire [31:0] grp_upzero_fu_442_bli_d0;
  reg [31:0] grp_upzero_fu_442_bli_q0;
  reg [31:0] zl1_i_reg_378;
  reg [2:0] dlt_pn_rec_i_reg_388;
  reg [31:0] zl1_i2_reg_399;
  reg [2:0] dlt_pn_rec_i2_reg_409;
  reg [4:0] ad_ptr_1_rec_reg_420;
  wire ap_CS_fsm_state29;
  reg [3:0] i_1_reg_431;
  reg grp_upzero_fu_442_ap_start_reg;
  wire [63:0] p_01_rec_i_cast_fu_545_p1;
  wire [63:0] tmp_s_fu_566_p1;
  wire [63:0] tmp_45_fu_576_p1;
  wire [63:0] tmp_i2_fu_762_p1;
  wire [63:0] p_01_rec_i2_cast_fu_1196_p1;
  wire [63:0] tmp_i6_fu_1384_p1;
  wire [63:0] ac_ptr_0_sum_cast_fu_1835_p1;
  wire [63:0] ad_ptr_0_sum7_cast_fu_1853_p1;
  wire signed [31:0] tmp_44_fu_686_p1;
  wire signed [31:0] tmp_64_cast_fu_860_p1;
  wire signed [31:0] tmp_51_fu_1403_p1;
  wire signed [31:0] tmp_70_cast_fu_1450_p1;
  wire signed [31:0] ih_assign_fu_529_p1;
  wire [31:0] nbl_assign_5_cast_fu_732_p1;
  wire [14:0] tmp_10_i_fu_840_p3;
  wire [31:0] dec_rlt_fu_874_p2;
  wire signed [31:0] apl2_assign_cast_fu_1118_p1;
  wire signed [31:0] apl1_12_cast_fu_1180_p1;
  wire [31:0] nbl_assign_6_cast_fu_1354_p1;
  wire [14:0] tmp_10_i2_fu_1430_p3;
  wire signed [31:0] apl2_assign_2_cast_fu_1720_p1;
  wire signed [31:0] apl1_16_cast_fu_1784_p1;
  wire [31:0] rh_fu_1801_p2;
  wire [0:0] exitcond_fu_1859_p2;
  wire [25:0] tmp_41_fu_519_p4;
  wire [3:0] tmp_1_cast_fu_557_p4;
  wire [31:0] tmp_72_fu_596_p2;
  wire [31:0] tmp_i7_fu_602_p2;
  wire signed [24:0] tmp_32_i_fu_608_p4;
  wire signed [12:0] wl_code_table_load_c_fu_622_p0;
  wire signed [12:0] tmp_13_fu_626_p0;
  wire signed [25:0] wd_cast_fu_618_p1;
  wire signed [25:0] wl_code_table_load_c_fu_622_p1;
  wire signed [24:0] tmp_13_fu_626_p1;
  wire [25:0] nbl_assign_4_fu_630_p2;
  wire signed [31:0] pl_fu_654_p0;
  wire signed [31:0] pl_fu_654_p1;
  wire signed [31:0] tmp_i1_fu_660_p0;
  wire signed [31:0] tmp_i1_fu_660_p1;
  wire signed [30:0] tmp_42_fu_1871_p2;
  wire signed [30:0] tmp_46_fu_1878_p2;
  wire [24:0] p_i_fu_708_p3;
  wire [0:0] tmp_18_i_fu_718_p2;
  wire [14:0] tmp_74_fu_714_p1;
  wire [14:0] nbl_assign_5_fu_724_p3;
  wire [4:0] wd1_fu_742_p4;
  wire [17:0] tmp_39_i_fu_767_p4;
  wire [31:0] tmp_i_31_fu_781_p2;
  wire [16:0] tmp_41_i_fu_785_p4;
  wire signed [18:0] tmp_20_i_cast_fu_795_p1;
  wire signed [18:0] tmp_i_cast_fu_777_p1;
  wire signed [18:0] dec_sl_fu_799_p2;
  wire signed [18:0] dl_cast_fu_816_p1;
  wire [3:0] tmp_9_i_fu_825_p2;
  wire [11:0] tmp_9_i_cast_cast_fu_830_p1;
  wire [11:0] wd3_fu_834_p2;
  wire signed [18:0] tmp_59_cast_fu_813_p1;
  wire [18:0] tmp_48_fu_854_p2;
  wire signed [31:0] dec_sl_cast_fu_805_p1;
  wire signed [31:0] tmp_i8_fu_904_p0;
  wire signed [31:0] tmp_i8_fu_904_p1;
  wire signed [31:0] tmp_5_i_fu_910_p0;
  wire signed [31:0] tmp_5_i_fu_910_p1;
  wire [31:0] wd2_fu_936_p2;
  wire [31:0] wd2_4_fu_949_p2;
  wire [0:0] tmp_76_fu_942_p3;
  wire [24:0] tmp_54_fu_965_p4;
  wire [24:0] tmp_53_fu_955_p4;
  wire [24:0] tmp_55_fu_975_p3;
  wire [0:0] tmp_77_fu_987_p3;
  wire [31:0] tmp_78_fu_1002_p2;
  wire [31:0] tmp_9_i4_fu_1008_p2;
  wire [24:0] tmp_19_i_fu_1014_p4;
  wire signed [25:0] wd2_15_cast_fu_983_p1;
  wire signed [25:0] tmp_1_i_cast_fu_1024_p1;
  wire [25:0] tmp4_fu_1028_p2;
  wire [26:0] tmp_8_i_cast_cast_fu_994_p3;
  wire signed [26:0] tmp4_cast_fu_1034_p1;
  wire [31:0] tmp_80_fu_1044_p2;
  wire [31:0] tmp_i9_fu_1050_p2;
  wire [0:0] tmp_2_i_fu_1066_p2;
  wire [26:0] p_i4_fu_1071_p3;
  wire [0:0] tmp_3_i_fu_1082_p2;
  wire [14:0] tmp_79_fu_1078_p1;
  wire signed [24:0] wd2_16_cast_fu_1096_p1;
  wire [24:0] tmp_4_i_cast_cast_fu_1099_p3;
  wire [24:0] tmp5_fu_1106_p2;
  wire [14:0] apl1_17_fu_1127_p2;
  wire [24:0] apl1_17_cast_fu_1136_p1;
  wire [0:0] tmp_6_i_fu_1140_p2;
  wire [24:0] wd3_0_apl1_i_fu_1145_p3;
  wire [15:0] apl1_17_cast1_fu_1132_p1;
  wire signed [24:0] apl1_11_cast_fu_1162_p1;
  wire [15:0] apl1_12_fu_1175_p3;
  wire [1:0] tmp_83_fu_1212_p1;
  wire [31:0] tmp_84_fu_1234_p2;
  wire [31:0] tmp_i2_35_fu_1240_p2;
  wire signed [24:0] tmp_36_i_fu_1246_p4;
  wire [31:0] tmp_15_fu_1260_p6;
  wire signed [31:0] wd_fu_1256_p1;
  wire signed [30:0] tmp_16_fu_1274_p1;
  wire [30:0] tmp_85_fu_1278_p1;
  wire [31:0] nbh_assign_2_fu_1282_p2;
  wire [14:0] tmp_49_fu_1315_p0;
  wire [31:0] tmp_49_fu_1315_p2;
  wire [30:0] p_i5_fu_1330_p3;
  wire [0:0] tmp_19_i3_fu_1340_p2;
  wire [14:0] tmp_87_fu_1336_p1;
  wire [14:0] nbl_assign_6_fu_1346_p3;
  wire [4:0] wd1_2_fu_1364_p4;
  wire [17:0] tmp_39_i2_fu_1389_p4;
  wire [3:0] tmp_9_i5_fu_1415_p2;
  wire [11:0] tmp_9_i5_cast_cast_fu_1420_p1;
  wire [11:0] wd3_5_fu_1424_p2;
  wire signed [18:0] tmp_69_cast_fu_1406_p1;
  wire [18:0] tmp_52_fu_1444_p2;
  wire signed [31:0] tmp_i3_fu_1472_p0;
  wire signed [31:0] tmp_i3_fu_1472_p1;
  wire signed [31:0] tmp_5_i5_fu_1478_p0;
  wire signed [31:0] tmp_5_i5_fu_1478_p1;
  wire [31:0] wd2_5_fu_1504_p2;
  wire [31:0] wd2_6_fu_1517_p2;
  wire [0:0] tmp_89_fu_1510_p3;
  wire [24:0] tmp_57_fu_1533_p4;
  wire [24:0] tmp_56_fu_1523_p4;
  wire [24:0] tmp_58_fu_1543_p3;
  wire [0:0] tmp_90_fu_1555_p3;
  wire [31:0] tmp_91_fu_1570_p2;
  wire [31:0] tmp_9_i6_fu_1576_p2;
  wire [24:0] tmp_19_i4_fu_1582_p4;
  wire signed [25:0] tmp_1_i2_cast_fu_1592_p1;
  wire signed [25:0] wd2_21_cast_fu_1551_p1;
  wire [25:0] tmp6_fu_1596_p2;
  wire signed [26:0] tmp6_cast_fu_1602_p1;
  wire [26:0] tmp_8_i2_cast_cast_fu_1562_p3;
  wire [31:0] tmp_93_fu_1612_p2;
  wire [31:0] tmp_i4_36_fu_1618_p2;
  wire signed [31:0] pl_2_fu_1638_p0;
  wire signed [31:0] pl_2_fu_1638_p1;
  wire signed [31:0] tmp_i4_fu_1644_p0;
  wire signed [31:0] tmp_i4_fu_1644_p1;
  wire [0:0] tmp_2_i2_fu_1650_p2;
  wire [26:0] p_i6_fu_1655_p3;
  wire [0:0] tmp_3_i2_fu_1666_p2;
  wire [14:0] tmp_92_fu_1662_p1;
  wire signed [24:0] wd2_22_cast_fu_1680_p1;
  wire [24:0] tmp7_fu_1690_p2;
  wire [24:0] tmp_4_i2_cast_cast_fu_1683_p3;
  wire [31:0] tmp_i1_34_fu_1702_p2;
  wire [16:0] tmp_41_i2_fu_1706_p4;
  wire [14:0] apl1_18_fu_1729_p2;
  wire [24:0] apl1_18_cast_fu_1738_p1;
  wire [0:0] tmp_6_i2_fu_1742_p2;
  wire [24:0] wd3_0_apl1_i2_fu_1747_p3;
  wire [15:0] apl1_18_cast9_fu_1734_p1;
  wire signed [24:0] apl1_15_cast_fu_1764_p1;
  wire signed [18:0] tmp_20_i5_cast_fu_1716_p1;
  wire [15:0] apl1_16_fu_1779_p3;
  wire signed [31:0] tmp8_cast_fu_1798_p1;
  wire [4:0] ac_ptr_0_sum_fu_1829_p2;
  wire [4:0] ad_ptr_0_sum7_fu_1847_p2;
  wire [14:0] tmp_42_fu_1871_p1;
  wire [30:0] extLd_cast_fu_670_p1;
  wire [14:0] tmp_46_fu_1878_p1;
  reg [28:0] ap_NS_fsm;
  wire [31:0] tmp_49_fu_1315_p00;
  wire [31:0] temp140;
  wire [31:0] temp142;
  wire [31:0] temp143;
  wire [31:0] temp144;
  wire [31:0] temp146;
  wire [31:0] temp147;
  wire [31:0] temp148;
  wire [31:0] temp150;
  wire [31:0] temp151;
  wire [31:0] temp152;
  wire [31:0] temp154;
  wire [31:0] temp155;
  wire [31:0] temp156;
  wire [31:0] temp158;
  wire [31:0] temp159;
  wire [31:0] temp160;
  wire [31:0] temp162;
  wire [31:0] temp163;
  wire [31:0] temp164;
  wire [31:0] temp166;
  wire [31:0] temp167;
  wire [31:0] temp168;
  wire [31:0] temp170;
  wire [31:0] temp171;
  wire [31:0] temp172;
  wire [31:0] temp174;
  wire [31:0] temp175;
  wire [31:0] temp176;
  wire [31:0] temp178;
  wire [31:0] temp179;
  input [109:0] working_key;

  initial begin
    #0 ap_CS_fsm = 29'd1;
    #0 dec_dlt = 32'd0;
    #0 dec_plt = 32'd0;
    #0 dec_dh = 32'd0;
    #0 dec_ph = 32'd0;
    #0 grp_upzero_fu_442_ap_start_reg = 1'b0;
  end


  encode_qq4_code4_dEe
  #(
    .DataWidth(16),
    .AddressRange(16),
    .AddressWidth(4)
  )
  qq4_code4_table_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(qq4_code4_table_address0),
    .ce0(qq4_code4_table_ce0),
    .q0(qq4_code4_table_q0)
  );


  decode_qq6_code6_kbM
  #(
    .DataWidth(16),
    .AddressRange(64),
    .AddressWidth(6)
  )
  qq6_code6_table_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(qq6_code6_table_address0),
    .ce0(qq6_code6_table_ce0),
    .q0(qq6_code6_table_q0)
  );


  encode_wl_code_taeOg
  #(
    .DataWidth(13),
    .AddressRange(16),
    .AddressWidth(4)
  )
  wl_code_table_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(wl_code_table_address0),
    .ce0(wl_code_table_ce0),
    .q0(wl_code_table_q0)
  );


  encode_ilb_table
  #(
    .DataWidth(12),
    .AddressRange(32),
    .AddressWidth(5)
  )
  ilb_table_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(ilb_table_address0),
    .ce0(ilb_table_ce0),
    .q0(ilb_table_q0)
  );


  upzero
  grp_upzero_fu_442
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_upzero_fu_442_ap_start),
    .ap_done(grp_upzero_fu_442_ap_done),
    .ap_idle(grp_upzero_fu_442_ap_idle),
    .ap_ready(grp_upzero_fu_442_ap_ready),
    .dlt(grp_upzero_fu_442_dlt),
    .dlti_address0(grp_upzero_fu_442_dlti_address0),
    .dlti_ce0(grp_upzero_fu_442_dlti_ce0),
    .dlti_we0(grp_upzero_fu_442_dlti_we0),
    .dlti_d0(grp_upzero_fu_442_dlti_d0),
    .dlti_q0(grp_upzero_fu_442_dlti_q0),
    .dlti_address1(grp_upzero_fu_442_dlti_address1),
    .dlti_ce1(grp_upzero_fu_442_dlti_ce1),
    .dlti_we1(grp_upzero_fu_442_dlti_we1),
    .dlti_d1(grp_upzero_fu_442_dlti_d1),
    .dlti_q1(grp_upzero_fu_442_dlti_q1),
    .bli_address0(grp_upzero_fu_442_bli_address0),
    .bli_ce0(grp_upzero_fu_442_bli_ce0),
    .bli_we0(grp_upzero_fu_442_bli_we0),
    .bli_d0(grp_upzero_fu_442_bli_d0),
    .bli_q0(grp_upzero_fu_442_bli_q0)
    .working_key(working_key)
  );


  adpcm_main_mux_42fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(32),
    .din1_WIDTH(32),
    .din2_WIDTH(32),
    .din3_WIDTH(32),
    .din4_WIDTH(2),
    .dout_WIDTH(32)
  )
  adpcm_main_mux_42fYi_U90
  (
    .din0(32'd4294959888),
    .din1(32'd4294965680),
    .din2(32'd7408),
    .din3(32'd1616),
    .din4(tmp_83_fu_1212_p1),
    .dout(tmp_14_fu_1216_p6)
  );


  adpcm_main_mux_42fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(32),
    .din1_WIDTH(32),
    .din2_WIDTH(32),
    .din3_WIDTH(32),
    .din4_WIDTH(2),
    .dout_WIDTH(32)
  )
  adpcm_main_mux_42fYi_U91
  (
    .din0(32'd798),
    .din1(32'd4294967082),
    .din2(32'd798),
    .din3(32'd4294967082),
    .din4(tmp_83_fu_1212_p1),
    .dout(tmp_15_fu_1260_p6)
  );


  adpcm_main_mul_mumb6
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(15),
    .dout_WIDTH(31)
  )
  adpcm_main_mul_mumb6_U92
  (
    .din0(qq4_code4_table_load_reg_1938),
    .din1(tmp_42_fu_1871_p1),
    .dout(tmp_42_fu_1871_p2)
  );


  adpcm_main_mul_mumb6
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(15),
    .dout_WIDTH(31)
  )
  adpcm_main_mul_mumb6_U93
  (
    .din0(qq6_code6_table_load_reg_1943),
    .din1(tmp_46_fu_1878_p1),
    .dout(tmp_46_fu_1878_p2)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_upzero_fu_442_ap_start_reg <= 1'b0;
    end else begin
      if((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state11)) begin
        grp_upzero_fu_442_ap_start_reg <= 1'b1;
      end else if(grp_upzero_fu_442_ap_ready == 1'b1) begin
        grp_upzero_fu_442_ap_start_reg <= 1'b0;
      end 
    end
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      if(working_key[41] == 1'b1) begin
        ad_ptr_1_rec_reg_420 <= 5'd0;
      end else begin
        ad_ptr_1_rec_reg_420 <= temp140;
      end
    end else if(1'b1 == ap_CS_fsm_state29) begin
      ad_ptr_1_rec_reg_420 <= p_rec_reg_2216;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state20) begin
      if(working_key[44] == 1'b1) begin
        dlt_pn_rec_i2_reg_409 <= temp144;
      end else begin
        dlt_pn_rec_i2_reg_409 <= p_01_rec_i2_reg_2063;
      end
    end else if(1'b1 == ap_CS_fsm_state16) begin
      dlt_pn_rec_i2_reg_409 <= 3'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state8) begin
      if(working_key[47] == 1'b1) begin
        dlt_pn_rec_i_reg_388 <= temp148;
      end else begin
        dlt_pn_rec_i_reg_388 <= p_01_rec_i_reg_1895;
      end
    end else if(1'b1 == ap_CS_fsm_state4) begin
      dlt_pn_rec_i_reg_388 <= 3'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      if(working_key[50] == 1'b1) begin
        i_1_reg_431 <= temp152;
      end else begin
        i_1_reg_431 <= 4'd0;
      end
    end else if(1'b1 == ap_CS_fsm_state29) begin
      i_1_reg_431 <= i_reg_2234;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state20) begin
      if(working_key[53] == 1'b1) begin
        zl1_i2_reg_399 <= zl_6_fu_1302_p2;
      end else begin
        zl1_i2_reg_399 <= temp156;
      end
    end else if(1'b1 == ap_CS_fsm_state16) begin
      zl1_i2_reg_399 <= zl_4_reg_2052;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state8) begin
      if(working_key[56] == 1'b1) begin
        zl1_i_reg_378 <= temp160;
      end else begin
        zl1_i_reg_378 <= zl_5_fu_587_p2;
      end
    end else if(1'b1 == ap_CS_fsm_state4) begin
      zl1_i_reg_378 <= zl_reg_1885;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state28) begin
      if(working_key[65] == 1'b1) begin
        accumc_addr_reg_2206 <= ac_ptr_0_sum_cast_fu_1835_p1;
        accumd_addr_reg_2211 <= ac_ptr_0_sum_cast_fu_1835_p1;
        i_reg_2234 <= i_fu_1865_p2;
        p_rec_reg_2216 <= p_rec_fu_1841_p2;
      end else begin
        accumc_addr_reg_2206 <= temp164;
        accumd_addr_reg_2211 <= temp168;
        i_reg_2234 <= temp172;
        p_rec_reg_2216 <= temp176;
      end
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state15) begin
      if(working_key[66] == 1'b1) begin
        apl1_11_reg_2042 <= apl1_11_fu_1156_p2;
        tmp_7_i_reg_2047 <= tmp_7_i_fu_1166_p2;
        tmp_82_reg_2037 <= tmp_82_fu_1152_p1;
        zl_4_reg_2052 <= grp_fu_493_p2;
      end else begin
        apl1_11_reg_2042 <= tmp_70_cast_fu_1450_p1;
        tmp_7_i_reg_2047 <= grp_upzero_fu_442_bli_we0;
        tmp_82_reg_2037 <= apl1_fu_1112_p2;
        zl_4_reg_2052 <= rl_cast_fu_1172_p1;
      end
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state25) begin
      if(working_key[67] == 1'b1) begin
        apl1_13_reg_2170 <= apl1_13_fu_1696_p2;
        apl2_assign_2_reg_2164 <= apl2_assign_2_fu_1672_p3;
        pl_2_reg_2154 <= pl_2_fu_1638_p2;
        tmp_i4_reg_2159 <= tmp_i4_fu_1644_p2;
      end else begin
        apl1_13_reg_2170 <= zl_4_reg_2052;
        apl2_assign_2_reg_2164 <= grp_fu_493_p2;
        pl_2_reg_2154 <= apl2_assign_fu_1088_p3;
        tmp_i4_reg_2159 <= grp_upzero_fu_442_dlti_address0;
      end
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state26) begin
      apl1_15_reg_2181 <= apl1_15_fu_1758_p2;
      tmp8_reg_2191 <= tmp8_fu_1774_p2;
      tmp_7_i2_reg_2186 <= tmp_7_i2_fu_1768_p2;
      tmp_95_reg_2176 <= tmp_95_fu_1754_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state14) begin
      apl1_reg_2031 <= apl1_fu_1112_p2;
      apl2_assign_reg_2025 <= apl2_assign_fu_1088_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state24) begin
      apl2_2_reg_2143 <= apl2_2_fu_1606_p2;
      tmp_21_i2_reg_2149 <= { { tmp_i4_36_fu_1618_p2[31:8] } };
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      apl2_reg_2014 <= apl2_fu_1038_p2;
      tmp_21_i_reg_2020 <= { { tmp_i9_fu_1050_p2[31:8] } };
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state22) begin
      dec_dh <= tmp_51_fu_1403_p1;
      dec_ph <= tmp_70_cast_fu_1450_p1;
      tmp_i19_cast_reg_2123 <= tmp_i19_cast_fu_1399_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state10) begin
      dec_dlt <= tmp_44_fu_686_p1;
      pl_reg_1958 <= pl_fu_654_p2;
      tmp_70_reg_1968 <= { { tmp_42_fu_1871_p2[30:15] } };
      tmp_71_reg_1974 <= { { tmp_46_fu_1878_p2[30:15] } };
      tmp_i1_reg_1963 <= tmp_i1_fu_660_p2;
      wd2_cast_reg_1979 <= { { nbl_assign_5_fu_724_p3[14:11] } };
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      dec_plt <= tmp_64_cast_fu_860_p1;
      rl_reg_1994 <= rl_fu_819_p2;
      tmp_43_reg_1989 <= tmp_43_fu_809_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond2_fu_1202_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state17)) begin
      nbh_assign_2_cast_reg_2086 <= nbh_assign_2_cast_fu_1288_p2;
      tmp_14_reg_2081 <= tmp_14_fu_1216_p6;
      tmp_86_reg_2091 <= nbh_assign_2_fu_1282_p2[32'd31];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      nbl_assign_4_cast_reg_1948 <= nbl_assign_4_cast_fu_636_p2;
      qq4_code4_table_load_reg_1938 <= qq4_code4_table_q0;
      qq6_code6_table_load_reg_1943 <= qq6_code6_table_q0;
      tmp_73_reg_1953 <= nbl_assign_4_fu_630_p2[32'd25];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state17) begin
      p_01_rec_i2_reg_2063 <= p_01_rec_i2_fu_1190_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      p_01_rec_i_reg_1895 <= p_01_rec_i_fu_539_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state2)) begin
      reg_477 <= dec_del_bpl_q0;
      reg_481 <= dec_del_dltx_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state14)) begin
      reg_485 <= dec_del_bph_q0;
      reg_489 <= dec_del_dhx_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      rl_cast_reg_2057 <= rl_cast_fu_1172_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state21) begin
      tmp_50_reg_2106 <= { { tmp_49_fu_1315_p2[31:15] } };
      wd2_17_cast_reg_2113 <= { { nbl_assign_6_fu_1346_p3[14:11] } };
    end 
  end


  always @(posedge ap_clk) begin
    if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state23)) begin
      tmp_5_i5_reg_2133 <= tmp_5_i5_fu_1478_p2;
      tmp_94_reg_2138 <= tmp_i3_fu_1472_p2[32'd31];
      tmp_i3_reg_2128 <= tmp_i3_fu_1472_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state12)) begin
      tmp_5_i_reg_2004 <= tmp_5_i_fu_910_p2;
      tmp_81_reg_2009 <= tmp_i8_fu_904_p2[32'd31];
      tmp_i8_reg_1999 <= tmp_i8_fu_904_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state19) begin
      tmp_i8_33_reg_2096 <= grp_fu_493_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      tmp_i_reg_1928 <= tmp_i_fu_581_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      xd_reg_2196 <= xd_fu_1819_p2;
      xs_reg_2201 <= xs_fu_1824_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      zl_reg_1885 <= zl_fu_499_p2;
    end 
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state29) begin
      accumc_address0 = accumc_addr_reg_2206;
    end else if((exitcond_fu_1859_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28)) begin
      accumc_address0 = 4'd0;
    end else if((exitcond_fu_1859_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state28)) begin
      accumc_address0 = ad_ptr_0_sum7_cast_fu_1853_p1;
    end else begin
      accumc_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state29) | (exitcond_fu_1859_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28) | (exitcond_fu_1859_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state28)) begin
      accumc_ce0 = 1'b1;
    end else begin
      accumc_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state29) begin
      accumc_d0 = accumc_q0;
    end else if((exitcond_fu_1859_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28)) begin
      accumc_d0 = xd_reg_2196;
    end else begin
      accumc_d0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state29) | (exitcond_fu_1859_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28)) begin
      accumc_we0 = 1'b1;
    end else begin
      accumc_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state29) begin
      accumd_address0 = accumd_addr_reg_2211;
    end else if((exitcond_fu_1859_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28)) begin
      accumd_address0 = 4'd0;
    end else if((exitcond_fu_1859_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state28)) begin
      accumd_address0 = ad_ptr_0_sum7_cast_fu_1853_p1;
    end else begin
      accumd_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state29) | (exitcond_fu_1859_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28) | (exitcond_fu_1859_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state28)) begin
      accumd_ce0 = 1'b1;
    end else begin
      accumd_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state29) begin
      accumd_d0 = accumd_q0;
    end else if((exitcond_fu_1859_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28)) begin
      accumd_d0 = xs_reg_2201;
    end else begin
      accumd_d0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state29) | (exitcond_fu_1859_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28)) begin
      accumd_we0 = 1'b1;
    end else begin
      accumd_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond_fu_1859_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28) | (ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond_fu_1859_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28)) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      dec_ah1_o = apl1_16_cast_fu_1784_p1;
    end else begin
      dec_ah1_o = dec_ah1_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      dec_ah1_o_ap_vld = 1'b1;
    end else begin
      dec_ah1_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state26) begin
      dec_ah2_o = apl2_assign_2_cast_fu_1720_p1;
    end else begin
      dec_ah2_o = dec_ah2_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state26) begin
      dec_ah2_o_ap_vld = 1'b1;
    end else begin
      dec_ah2_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      dec_al1_o = apl1_12_cast_fu_1180_p1;
    end else begin
      dec_al1_o = dec_al1_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      dec_al1_o_ap_vld = 1'b1;
    end else begin
      dec_al1_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state15) begin
      dec_al2_o = apl2_assign_cast_fu_1118_p1;
    end else begin
      dec_al2_o = dec_al2_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state15) begin
      dec_al2_o_ap_vld = 1'b1;
    end else begin
      dec_al2_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state17) begin
      dec_del_bph_address0 = p_01_rec_i2_cast_fu_1196_p1;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      dec_del_bph_address0 = 3'd0;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      dec_del_bph_address0 = grp_upzero_fu_442_bli_address0;
    end else begin
      dec_del_bph_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state13)) begin
      dec_del_bph_ce0 = 1'b1;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      dec_del_bph_ce0 = grp_upzero_fu_442_bli_ce0;
    end else begin
      dec_del_bph_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state23) begin
      dec_del_bph_we0 = grp_upzero_fu_442_bli_we0;
    end else begin
      dec_del_bph_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      dec_del_bpl_address0 = p_01_rec_i_cast_fu_545_p1;
    end else if(1'b1 == ap_CS_fsm_state1) begin
      dec_del_bpl_address0 = 3'd0;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      dec_del_bpl_address0 = grp_upzero_fu_442_bli_address0;
    end else begin
      dec_del_bpl_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state5) | (ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      dec_del_bpl_ce0 = 1'b1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      dec_del_bpl_ce0 = grp_upzero_fu_442_bli_ce0;
    end else begin
      dec_del_bpl_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      dec_del_bpl_we0 = grp_upzero_fu_442_bli_we0;
    end else begin
      dec_del_bpl_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state17) begin
      dec_del_dhx_address0 = p_01_rec_i2_cast_fu_1196_p1;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      dec_del_dhx_address0 = 3'd0;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      dec_del_dhx_address0 = grp_upzero_fu_442_dlti_address0;
    end else begin
      dec_del_dhx_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state13)) begin
      dec_del_dhx_ce0 = 1'b1;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      dec_del_dhx_ce0 = grp_upzero_fu_442_dlti_ce0;
    end else begin
      dec_del_dhx_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state23) begin
      dec_del_dhx_ce1 = grp_upzero_fu_442_dlti_ce1;
    end else begin
      dec_del_dhx_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state23) begin
      dec_del_dhx_we0 = grp_upzero_fu_442_dlti_we0;
    end else begin
      dec_del_dhx_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state23) begin
      dec_del_dhx_we1 = grp_upzero_fu_442_dlti_we1;
    end else begin
      dec_del_dhx_we1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      dec_del_dltx_address0 = p_01_rec_i_cast_fu_545_p1;
    end else if(1'b1 == ap_CS_fsm_state1) begin
      dec_del_dltx_address0 = 3'd0;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      dec_del_dltx_address0 = grp_upzero_fu_442_dlti_address0;
    end else begin
      dec_del_dltx_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state5) | (ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      dec_del_dltx_ce0 = 1'b1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      dec_del_dltx_ce0 = grp_upzero_fu_442_dlti_ce0;
    end else begin
      dec_del_dltx_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      dec_del_dltx_ce1 = grp_upzero_fu_442_dlti_ce1;
    end else begin
      dec_del_dltx_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      dec_del_dltx_we0 = grp_upzero_fu_442_dlti_we0;
    end else begin
      dec_del_dltx_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      dec_del_dltx_we1 = grp_upzero_fu_442_dlti_we1;
    end else begin
      dec_del_dltx_we1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state22) begin
      dec_deth_o = tmp_10_i2_fu_1430_p3;
    end else begin
      dec_deth_o = dec_deth_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state22) begin
      dec_deth_o_ap_vld = 1'b1;
    end else begin
      dec_deth_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      dec_detl_o = tmp_10_i_fu_840_p3;
    end else begin
      dec_detl_o = dec_detl_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      dec_detl_o_ap_vld = 1'b1;
    end else begin
      dec_detl_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state21) begin
      dec_nbh_o = nbl_assign_6_cast_fu_1354_p1;
    end else begin
      dec_nbh_o = dec_nbh_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state21) begin
      dec_nbh_o_ap_vld = 1'b1;
    end else begin
      dec_nbh_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state10) begin
      dec_nbl_o = nbl_assign_5_cast_fu_732_p1;
    end else begin
      dec_nbl_o = dec_nbl_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state10) begin
      dec_nbl_o_ap_vld = 1'b1;
    end else begin
      dec_nbl_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state23)) begin
      dec_ph1_o = dec_ph;
    end else begin
      dec_ph1_o = dec_ph1_i;
    end
  end


  always @(*) begin
    if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state23)) begin
      dec_ph1_o_ap_vld = 1'b1;
    end else begin
      dec_ph1_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state23)) begin
      dec_ph2_o = dec_ph1_i;
    end else begin
      dec_ph2_o = dec_ph2_i;
    end
  end


  always @(*) begin
    if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state23)) begin
      dec_ph2_o_ap_vld = 1'b1;
    end else begin
      dec_ph2_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state12)) begin
      dec_plt1_o = dec_plt;
    end else begin
      dec_plt1_o = dec_plt1_i;
    end
  end


  always @(*) begin
    if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state12)) begin
      dec_plt1_o_ap_vld = 1'b1;
    end else begin
      dec_plt1_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state12)) begin
      dec_plt2_o = dec_plt1_i;
    end else begin
      dec_plt2_o = dec_plt2_i;
    end
  end


  always @(*) begin
    if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state12)) begin
      dec_plt2_o_ap_vld = 1'b1;
    end else begin
      dec_plt2_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      dec_rh1_o = rh_fu_1801_p2;
    end else begin
      dec_rh1_o = dec_rh1_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      dec_rh1_o_ap_vld = 1'b1;
    end else begin
      dec_rh1_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      dec_rh2_o = dec_rh1_i;
    end else begin
      dec_rh2_o = dec_rh2_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      dec_rh2_o_ap_vld = 1'b1;
    end else begin
      dec_rh2_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      dec_rlt1_o = dec_rlt_fu_874_p2;
    end else begin
      dec_rlt1_o = dec_rlt1_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      dec_rlt1_o_ap_vld = 1'b1;
    end else begin
      dec_rlt1_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      dec_rlt2_o = dec_rlt1_i;
    end else begin
      dec_rlt2_o = dec_rlt2_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      dec_rlt2_o_ap_vld = 1'b1;
    end else begin
      dec_rlt2_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state23) begin
      grp_upzero_fu_442_bli_q0 = dec_del_bph_q0;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      grp_upzero_fu_442_bli_q0 = dec_del_bpl_q0;
    end else begin
      grp_upzero_fu_442_bli_q0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state23) begin
      grp_upzero_fu_442_dlt = tmp_50_reg_2106;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      grp_upzero_fu_442_dlt = tmp_43_reg_1989;
    end else begin
      grp_upzero_fu_442_dlt = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state23) begin
      grp_upzero_fu_442_dlti_q0 = dec_del_dhx_q0;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      grp_upzero_fu_442_dlti_q0 = dec_del_dltx_q0;
    end else begin
      grp_upzero_fu_442_dlti_q0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state23) begin
      grp_upzero_fu_442_dlti_q1 = dec_del_dhx_q1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      grp_upzero_fu_442_dlti_q1 = dec_del_dltx_q1;
    end else begin
      grp_upzero_fu_442_dlti_q1 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state4) begin
      ih_o = ih_assign_fu_529_p1;
    end else begin
      ih_o = ih_i;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state4) begin
      ih_o_ap_vld = 1'b1;
    end else begin
      ih_o_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state21) begin
      ilb_table_address0 = tmp_i6_fu_1384_p1;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      ilb_table_address0 = tmp_i2_fu_762_p1;
    end else begin
      ilb_table_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state10)) begin
      ilb_table_ce0 = 1'b1;
    end else begin
      ilb_table_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      qq4_code4_table_ce0 = 1'b1;
    end else begin
      qq4_code4_table_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      qq6_code6_table_ce0 = 1'b1;
    end else begin
      qq6_code6_table_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      wl_code_table_ce0 = 1'b1;
    end else begin
      wl_code_table_ce0 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        ap_NS_fsm = ap_ST_fsm_state3;
      end
      ap_ST_fsm_state3: begin
        ap_NS_fsm = ap_ST_fsm_state4;
      end
      ap_ST_fsm_state4: begin
        ap_NS_fsm = ap_ST_fsm_state5;
      end
      ap_ST_fsm_state5: begin
        if((exitcond3_fu_551_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state5)) begin
          ap_NS_fsm = ap_ST_fsm_state9;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end
      end
      ap_ST_fsm_state6: begin
        ap_NS_fsm = ap_ST_fsm_state7;
      end
      ap_ST_fsm_state7: begin
        ap_NS_fsm = ap_ST_fsm_state8;
      end
      ap_ST_fsm_state8: begin
        ap_NS_fsm = ap_ST_fsm_state5;
      end
      ap_ST_fsm_state9: begin
        ap_NS_fsm = ap_ST_fsm_state10;
      end
      ap_ST_fsm_state10: begin
        ap_NS_fsm = ap_ST_fsm_state11;
      end
      ap_ST_fsm_state11: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      ap_ST_fsm_state12: begin
        if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state12)) begin
          ap_NS_fsm = ap_ST_fsm_state13;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state12;
        end
      end
      ap_ST_fsm_state13: begin
        ap_NS_fsm = ap_ST_fsm_state14;
      end
      ap_ST_fsm_state14: begin
        ap_NS_fsm = ap_ST_fsm_state15;
      end
      ap_ST_fsm_state15: begin
        ap_NS_fsm = ap_ST_fsm_state16;
      end
      ap_ST_fsm_state16: begin
        ap_NS_fsm = ap_ST_fsm_state17;
      end
      ap_ST_fsm_state17: begin
        if((exitcond2_fu_1202_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state17)) begin
          ap_NS_fsm = ap_ST_fsm_state21;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state18;
        end
      end
      ap_ST_fsm_state18: begin
        ap_NS_fsm = ap_ST_fsm_state19;
      end
      ap_ST_fsm_state19: begin
        ap_NS_fsm = ap_ST_fsm_state20;
      end
      ap_ST_fsm_state20: begin
        ap_NS_fsm = ap_ST_fsm_state17;
      end
      ap_ST_fsm_state21: begin
        ap_NS_fsm = ap_ST_fsm_state22;
      end
      ap_ST_fsm_state22: begin
        ap_NS_fsm = ap_ST_fsm_state23;
      end
      ap_ST_fsm_state23: begin
        if((grp_upzero_fu_442_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state23)) begin
          ap_NS_fsm = ap_ST_fsm_state24;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state23;
        end
      end
      ap_ST_fsm_state24: begin
        ap_NS_fsm = ap_ST_fsm_state25;
      end
      ap_ST_fsm_state25: begin
        ap_NS_fsm = ap_ST_fsm_state26;
      end
      ap_ST_fsm_state26: begin
        ap_NS_fsm = ap_ST_fsm_state27;
      end
      ap_ST_fsm_state27: begin
        ap_NS_fsm = ap_ST_fsm_state28;
      end
      ap_ST_fsm_state28: begin
        if((exitcond_fu_1859_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28)) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state29;
        end
      end
      ap_ST_fsm_state29: begin
        ap_NS_fsm = ap_ST_fsm_state28;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign ac_ptr_0_sum_cast_fu_1835_p1 = ac_ptr_0_sum_fu_1829_p2;
  assign ac_ptr_0_sum_fu_1829_p2 = ad_ptr_1_rec_reg_420 + 5'd10;
  assign ad_ptr_0_sum7_cast_fu_1853_p1 = ad_ptr_0_sum7_fu_1847_p2;
  assign ad_ptr_0_sum7_fu_1847_p2 = ad_ptr_1_rec_reg_420 + 5'd9;
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];
  assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];
  assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];
  assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];
  assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];
  assign ap_CS_fsm_state21 = ap_CS_fsm[32'd20];
  assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];
  assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];
  assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];
  assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];
  assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];
  assign ap_CS_fsm_state27 = ap_CS_fsm[32'd26];
  assign ap_CS_fsm_state28 = ap_CS_fsm[32'd27];
  assign ap_CS_fsm_state29 = ap_CS_fsm[32'd28];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign apl1_11_cast_fu_1162_p1 = apl1_11_fu_1156_p2;
  assign apl1_11_fu_1156_p2 = 16'd0 - apl1_17_cast1_fu_1132_p1;
  assign apl1_12_cast_fu_1180_p1 = $signed(apl1_12_fu_1175_p3);
  assign apl1_12_fu_1175_p3 = (tmp_7_i_reg_2047[0:0] === 1'b1)? apl1_11_reg_2042 : tmp_82_reg_2037;
  assign apl1_13_fu_1696_p2 = tmp7_fu_1690_p2 + tmp_4_i2_cast_cast_fu_1683_p3;
  assign apl1_15_cast_fu_1764_p1 = apl1_15_fu_1758_p2;
  assign apl1_15_fu_1758_p2 = 16'd0 - apl1_18_cast9_fu_1734_p1;
  assign apl1_16_cast_fu_1784_p1 = $signed(apl1_16_fu_1779_p3);
  assign apl1_16_fu_1779_p3 = (tmp_7_i2_reg_2186[0:0] === 1'b1)? apl1_15_reg_2181 : tmp_95_reg_2176;
  assign apl1_17_cast1_fu_1132_p1 = apl1_17_fu_1127_p2;
  assign apl1_17_cast_fu_1136_p1 = apl1_17_fu_1127_p2;
  assign apl1_17_fu_1127_p2 = $signed(15'd15360) - $signed(apl2_assign_reg_2025);
  assign apl1_18_cast9_fu_1734_p1 = apl1_18_fu_1729_p2;
  assign apl1_18_cast_fu_1738_p1 = apl1_18_fu_1729_p2;
  assign apl1_18_fu_1729_p2 = $signed(15'd15360) - $signed(apl2_assign_2_reg_2164);
  assign apl1_fu_1112_p2 = tmp_4_i_cast_cast_fu_1099_p3 + tmp5_fu_1106_p2;
  assign apl2_2_fu_1606_p2 = $signed(tmp6_cast_fu_1602_p1) + $signed(tmp_8_i2_cast_cast_fu_1562_p3);
  assign apl2_assign_2_cast_fu_1720_p1 = apl2_assign_2_reg_2164;
  assign apl2_assign_2_fu_1672_p3 = (tmp_3_i2_fu_1666_p2[0:0] === 1'b1)? 15'd20480 : tmp_92_fu_1662_p1;
  assign apl2_assign_cast_fu_1118_p1 = apl2_assign_reg_2025;
  assign apl2_assign_fu_1088_p3 = (tmp_3_i_fu_1082_p2[0:0] === 1'b1)? 15'd20480 : tmp_79_fu_1078_p1;
  assign apl2_fu_1038_p2 = $signed(tmp_8_i_cast_cast_fu_994_p3) + $signed(tmp4_cast_fu_1034_p1);
  assign dec_del_bph_d0 = grp_upzero_fu_442_bli_d0;
  assign dec_del_bpl_d0 = grp_upzero_fu_442_bli_d0;
  assign dec_del_dhx_address1 = grp_upzero_fu_442_dlti_address1;
  assign dec_del_dhx_d0 = grp_upzero_fu_442_dlti_d0;
  assign dec_del_dhx_d1 = grp_upzero_fu_442_dlti_d1;
  assign dec_del_dltx_address1 = grp_upzero_fu_442_dlti_address1;
  assign dec_del_dltx_d0 = grp_upzero_fu_442_dlti_d0;
  assign dec_del_dltx_d1 = grp_upzero_fu_442_dlti_d1;
  assign dec_rlt_fu_874_p2 = $signed(dec_sl_cast_fu_805_p1) + $signed(dec_dlt);
  assign dec_sl_cast_fu_805_p1 = dec_sl_fu_799_p2;
  assign dec_sl_fu_799_p2 = $signed(tmp_20_i_cast_fu_795_p1) + $signed(tmp_i_cast_fu_777_p1);
  assign dl_cast_fu_816_p1 = $signed(tmp_71_reg_1974);
  assign exitcond2_fu_1202_p2 = (dlt_pn_rec_i2_reg_409 == 3'd5)? 1'b1 : 1'b0;
  assign exitcond3_fu_551_p2 = (dlt_pn_rec_i_reg_388 == 3'd5)? 1'b1 : 1'b0;
  assign exitcond_fu_1859_p2 = (i_1_reg_431 == 4'd10)? 1'b1 : 1'b0;
  assign extLd_cast_fu_670_p1 = dec_detl_i;
  assign grp_fu_493_p2 = $signed(reg_489) * $signed(reg_485);
  assign grp_upzero_fu_442_ap_start = grp_upzero_fu_442_ap_start_reg;
  assign i_fu_1865_p2 = i_1_reg_431 + 4'd1;
  assign ih_assign_fu_529_p1 = $signed(tmp_41_fu_519_p4);
  assign nbh_assign_2_cast_fu_1288_p2 = $signed(tmp_16_fu_1274_p1) + $signed(tmp_85_fu_1278_p1);
  assign nbh_assign_2_fu_1282_p2 = $signed(tmp_15_fu_1260_p6) + $signed(wd_fu_1256_p1);
  assign nbl_assign_4_cast_fu_636_p2 = $signed(tmp_13_fu_626_p1) + $signed(tmp_32_i_fu_608_p4);
  assign nbl_assign_4_fu_630_p2 = $signed(wd_cast_fu_618_p1) + $signed(wl_code_table_load_c_fu_622_p1);
  assign nbl_assign_5_cast_fu_732_p1 = nbl_assign_5_fu_724_p3;
  assign nbl_assign_5_fu_724_p3 = (tmp_18_i_fu_718_p2[0:0] === 1'b1)? 15'd18432 : tmp_74_fu_714_p1;
  assign nbl_assign_6_cast_fu_1354_p1 = nbl_assign_6_fu_1346_p3;
  assign nbl_assign_6_fu_1346_p3 = (tmp_19_i3_fu_1340_p2[0:0] === 1'b1)? 15'd22528 : tmp_87_fu_1336_p1;
  assign p_01_rec_i2_cast_fu_1196_p1 = p_01_rec_i2_fu_1190_p2;
  assign p_01_rec_i2_fu_1190_p2 = dlt_pn_rec_i2_reg_409 + 3'd1;
  assign p_01_rec_i_cast_fu_545_p1 = p_01_rec_i_fu_539_p2;
  assign p_01_rec_i_fu_539_p2 = dlt_pn_rec_i_reg_388 + 3'd1;
  assign p_i4_fu_1071_p3 = (tmp_2_i_fu_1066_p2[0:0] === 1'b1)? 27'd12288 : apl2_reg_2014;
  assign p_i5_fu_1330_p3 = (tmp_86_reg_2091[0:0] === 1'b1)? 31'd0 : nbh_assign_2_cast_reg_2086;
  assign p_i6_fu_1655_p3 = (tmp_2_i2_fu_1650_p2[0:0] === 1'b1)? 27'd12288 : apl2_2_reg_2143;
  assign p_i_fu_708_p3 = (tmp_73_reg_1953[0:0] === 1'b1)? 25'd0 : nbl_assign_4_cast_reg_1948;
  assign p_rec_fu_1841_p2 = $signed(ad_ptr_1_rec_reg_420) + $signed(5'd31);
  assign pl_2_fu_1638_p0 = dec_ah1_i;
  assign pl_2_fu_1638_p1 = dec_rh1_i;
  assign pl_2_fu_1638_p2 = $signed(pl_2_fu_1638_p0) * $signed(pl_2_fu_1638_p1);
  assign pl_fu_654_p0 = dec_rlt1_i;
  assign pl_fu_654_p1 = dec_al1_i;
  assign pl_fu_654_p2 = $signed(pl_fu_654_p0) * $signed(pl_fu_654_p1);
  assign qq4_code4_table_address0 = tmp_s_fu_566_p1;
  assign qq6_code6_table_address0 = tmp_45_fu_576_p1;
  assign rh_fu_1801_p2 = $signed(tmp8_cast_fu_1798_p1) + $signed(dec_dh);
  assign rl_cast_fu_1172_p1 = $signed(rl_reg_1994);
  assign rl_fu_819_p2 = $signed(dl_cast_fu_816_p1) + $signed(dec_sl_fu_799_p2);
  assign tmp4_cast_fu_1034_p1 = $signed(tmp4_fu_1028_p2);
  assign tmp4_fu_1028_p2 = $signed(wd2_15_cast_fu_983_p1) + $signed(tmp_1_i_cast_fu_1024_p1);
  assign tmp5_fu_1106_p2 = $signed(25'd192) + $signed(wd2_16_cast_fu_1096_p1);
  assign tmp6_cast_fu_1602_p1 = $signed(tmp6_fu_1596_p2);
  assign tmp6_fu_1596_p2 = $signed(tmp_1_i2_cast_fu_1592_p1) + $signed(wd2_21_cast_fu_1551_p1);
  assign tmp7_fu_1690_p2 = $signed(25'd192) + $signed(wd2_22_cast_fu_1680_p1);
  assign tmp8_cast_fu_1798_p1 = $signed(tmp8_reg_2191);
  assign tmp8_fu_1774_p2 = $signed(tmp_i19_cast_reg_2123) + $signed(tmp_20_i5_cast_fu_1716_p1);
  assign tmp_10_i2_fu_1430_p3 = { { wd3_5_fu_1424_p2 }, { 3'd0 } };
  assign tmp_10_i_fu_840_p3 = { { wd3_fu_834_p2 }, { 3'd0 } };
  assign tmp_13_fu_626_p0 = wl_code_table_q0;
  assign tmp_13_fu_626_p1 = tmp_13_fu_626_p0;
  assign tmp_16_fu_1274_p1 = tmp_36_i_fu_1246_p4;
  assign tmp_18_i_fu_718_p2 = (p_i_fu_708_p3 > 25'd18432)? 1'b1 : 1'b0;
  assign tmp_19_i3_fu_1340_p2 = (p_i5_fu_1330_p3 > 31'd22528)? 1'b1 : 1'b0;
  assign tmp_19_i4_fu_1582_p4 = { { tmp_9_i6_fu_1576_p2[31:7] } };
  assign tmp_19_i_fu_1014_p4 = { { tmp_9_i4_fu_1008_p2[31:7] } };
  assign tmp_1_cast_fu_557_p4 = { { input_r[5:2] } };
  assign tmp_1_i2_cast_fu_1592_p1 = $signed(tmp_19_i4_fu_1582_p4);
  assign tmp_1_i_cast_fu_1024_p1 = $signed(tmp_19_i_fu_1014_p4);
  assign tmp_20_i5_cast_fu_1716_p1 = $signed(tmp_41_i2_fu_1706_p4);
  assign tmp_20_i_cast_fu_795_p1 = $signed(tmp_41_i_fu_785_p4);
  assign tmp_2_i2_fu_1650_p2 = ($signed(apl2_2_reg_2143) > $signed(27'd12288))? 1'b1 : 1'b0;
  assign tmp_2_i_fu_1066_p2 = ($signed(apl2_reg_2014) > $signed(27'd12288))? 1'b1 : 1'b0;
  assign tmp_32_i_fu_608_p4 = { { tmp_i7_fu_602_p2[31:7] } };
  assign tmp_36_i_fu_1246_p4 = { { tmp_i2_35_fu_1240_p2[31:7] } };
  assign tmp_39_i2_fu_1389_p4 = { { zl1_i2_reg_399[31:14] } };
  assign tmp_39_i_fu_767_p4 = { { zl1_i_reg_378[31:14] } };
  assign tmp_3_i2_fu_1666_p2 = ($signed(p_i6_fu_1655_p3) < $signed(27'd134205440))? 1'b1 : 1'b0;
  assign tmp_3_i_fu_1082_p2 = ($signed(p_i4_fu_1071_p3) < $signed(27'd134205440))? 1'b1 : 1'b0;
  assign tmp_41_fu_519_p4 = { { input_r[31:6] } };
  assign tmp_41_i2_fu_1706_p4 = { { tmp_i1_34_fu_1702_p2[30:14] } };
  assign tmp_41_i_fu_785_p4 = { { tmp_i_31_fu_781_p2[30:14] } };
  assign tmp_42_fu_1871_p1 = extLd_cast_fu_670_p1;
  assign tmp_43_fu_809_p1 = tmp_70_reg_1968;
  assign tmp_44_fu_686_p1 = tmp_70_fu_677_p4;
  assign tmp_45_fu_576_p1 = il;
  assign tmp_46_fu_1878_p1 = extLd_cast_fu_670_p1;
  assign tmp_48_fu_854_p2 = $signed(tmp_59_cast_fu_813_p1) + $signed(tmp_i_cast_fu_777_p1);
  assign tmp_49_fu_1315_p0 = tmp_49_fu_1315_p00;
  assign tmp_49_fu_1315_p00 = dec_deth_i;
  assign tmp_49_fu_1315_p2 = $signed({ { 1'b0 }, { tmp_49_fu_1315_p0 } }) * $signed(tmp_14_reg_2081);
  assign tmp_4_i2_cast_cast_fu_1683_p3 = (tmp_94_reg_2138[0:0] === 1'b1)? 25'd33554048 : 25'd0;
  assign tmp_4_i_cast_cast_fu_1099_p3 = (tmp_81_reg_2009[0:0] === 1'b1)? 25'd33554048 : 25'd0;
  assign tmp_51_fu_1403_p1 = tmp_50_reg_2106;
  assign tmp_52_fu_1444_p2 = $signed(tmp_i19_cast_fu_1399_p1) + $signed(tmp_69_cast_fu_1406_p1);
  assign tmp_53_fu_955_p4 = { { wd2_4_fu_949_p2[31:7] } };
  assign tmp_54_fu_965_p4 = { { dec_al1_i[29:5] } };
  assign tmp_55_fu_975_p3 = (tmp_76_fu_942_p3[0:0] === 1'b1)? tmp_54_fu_965_p4 : tmp_53_fu_955_p4;
  assign tmp_56_fu_1523_p4 = { { wd2_6_fu_1517_p2[31:7] } };
  assign tmp_57_fu_1533_p4 = { { dec_ah1_i[29:5] } };
  assign tmp_58_fu_1543_p3 = (tmp_89_fu_1510_p3[0:0] === 1'b1)? tmp_57_fu_1533_p4 : tmp_56_fu_1523_p4;
  assign tmp_59_cast_fu_813_p1 = tmp_70_reg_1968;
  assign tmp_5_i5_fu_1478_p0 = dec_ph;
  assign tmp_5_i5_fu_1478_p1 = dec_ph2_i;
  assign tmp_5_i5_fu_1478_p2 = $signed(tmp_5_i5_fu_1478_p0) * $signed(tmp_5_i5_fu_1478_p1);
  assign tmp_5_i_fu_910_p0 = dec_plt2_i;
  assign tmp_5_i_fu_910_p1 = dec_plt;
  assign tmp_5_i_fu_910_p2 = $signed(tmp_5_i_fu_910_p0) * $signed(tmp_5_i_fu_910_p1);
  assign tmp_64_cast_fu_860_p1 = $signed(tmp_48_fu_854_p2);
  assign tmp_69_cast_fu_1406_p1 = tmp_50_reg_2106;
  assign tmp_6_i2_fu_1742_p2 = ($signed(apl1_13_reg_2170) > $signed(apl1_18_cast_fu_1738_p1))? 1'b1 : 1'b0;
  assign tmp_6_i_fu_1140_p2 = ($signed(apl1_reg_2031) > $signed(apl1_17_cast_fu_1136_p1))? 1'b1 : 1'b0;
  assign tmp_70_cast_fu_1450_p1 = $signed(tmp_52_fu_1444_p2);
  assign tmp_70_fu_677_p4 = { { tmp_42_fu_1871_p2[30:15] } };
  assign tmp_72_fu_596_p2 = dec_nbl_i << 32'd7;
  assign tmp_74_fu_714_p1 = p_i_fu_708_p3[14:0];
  assign tmp_76_fu_942_p3 = tmp_i8_reg_1999[32'd31];
  assign tmp_77_fu_987_p3 = tmp_5_i_reg_2004[32'd31];
  assign tmp_78_fu_1002_p2 = dec_al2_i << 32'd7;
  assign tmp_79_fu_1078_p1 = p_i4_fu_1071_p3[14:0];
  assign tmp_7_i2_fu_1768_p2 = ($signed(wd3_0_apl1_i2_fu_1747_p3) < $signed(apl1_15_cast_fu_1764_p1))? 1'b1 : 1'b0;
  assign tmp_7_i_fu_1166_p2 = ($signed(wd3_0_apl1_i_fu_1145_p3) < $signed(apl1_11_cast_fu_1162_p1))? 1'b1 : 1'b0;
  assign tmp_80_fu_1044_p2 = dec_al1_i << 32'd8;
  assign tmp_82_fu_1152_p1 = wd3_0_apl1_i_fu_1145_p3[15:0];
  assign tmp_83_fu_1212_p1 = ih_i[1:0];
  assign tmp_84_fu_1234_p2 = dec_nbh_i << 32'd7;
  assign tmp_85_fu_1278_p1 = tmp_15_fu_1260_p6[30:0];
  assign tmp_87_fu_1336_p1 = p_i5_fu_1330_p3[14:0];
  assign tmp_89_fu_1510_p3 = tmp_i3_reg_2128[32'd31];
  assign tmp_8_i2_cast_cast_fu_1562_p3 = (tmp_90_fu_1555_p3[0:0] === 1'b1)? 27'd134217600 : 27'd128;
  assign tmp_8_i_cast_cast_fu_994_p3 = (tmp_77_fu_987_p3[0:0] === 1'b1)? 27'd134217600 : 27'd128;
  assign tmp_90_fu_1555_p3 = tmp_5_i5_reg_2133[32'd31];
  assign tmp_91_fu_1570_p2 = dec_ah2_i << 32'd7;
  assign tmp_92_fu_1662_p1 = p_i6_fu_1655_p3[14:0];
  assign tmp_93_fu_1612_p2 = dec_ah1_i << 32'd8;
  assign tmp_95_fu_1754_p1 = wd3_0_apl1_i2_fu_1747_p3[15:0];
  assign tmp_9_i4_fu_1008_p2 = tmp_78_fu_1002_p2 - dec_al2_i;
  assign tmp_9_i5_cast_cast_fu_1420_p1 = tmp_9_i5_fu_1415_p2;
  assign tmp_9_i5_fu_1415_p2 = $signed(4'd11) - $signed(wd2_17_cast_reg_2113);
  assign tmp_9_i6_fu_1576_p2 = tmp_91_fu_1570_p2 - dec_ah2_i;
  assign tmp_9_i_cast_cast_fu_830_p1 = tmp_9_i_fu_825_p2;
  assign tmp_9_i_fu_825_p2 = $signed(4'd9) - $signed(wd2_cast_reg_1979);
  assign tmp_i19_cast_fu_1399_p1 = $signed(tmp_39_i2_fu_1389_p4);
  assign tmp_i1_34_fu_1702_p2 = tmp_i4_reg_2159 + pl_2_reg_2154;
  assign tmp_i1_fu_660_p0 = dec_rlt2_i;
  assign tmp_i1_fu_660_p1 = dec_al2_i;
  assign tmp_i1_fu_660_p2 = $signed(tmp_i1_fu_660_p0) * $signed(tmp_i1_fu_660_p1);
  assign tmp_i2_35_fu_1240_p2 = tmp_84_fu_1234_p2 - dec_nbh_i;
  assign tmp_i2_fu_762_p1 = wd1_fu_742_p4;
  assign tmp_i3_fu_1472_p0 = dec_ph;
  assign tmp_i3_fu_1472_p1 = dec_ph1_i;
  assign tmp_i3_fu_1472_p2 = $signed(tmp_i3_fu_1472_p0) * $signed(tmp_i3_fu_1472_p1);
  assign tmp_i4_36_fu_1618_p2 = tmp_93_fu_1612_p2 - dec_ah1_i;
  assign tmp_i4_fu_1644_p0 = dec_ah2_i;
  assign tmp_i4_fu_1644_p1 = dec_rh2_i;
  assign tmp_i4_fu_1644_p2 = $signed(tmp_i4_fu_1644_p0) * $signed(tmp_i4_fu_1644_p1);
  assign tmp_i6_fu_1384_p1 = wd1_2_fu_1364_p4;
  assign tmp_i7_fu_602_p2 = tmp_72_fu_596_p2 - dec_nbl_i;
  assign tmp_i8_fu_904_p0 = dec_plt1_i;
  assign tmp_i8_fu_904_p1 = dec_plt;
  assign tmp_i8_fu_904_p2 = $signed(tmp_i8_fu_904_p0) * $signed(tmp_i8_fu_904_p1);
  assign tmp_i9_fu_1050_p2 = tmp_80_fu_1044_p2 - dec_al1_i;
  assign tmp_i_31_fu_781_p2 = pl_reg_1958 + tmp_i1_reg_1963;
  assign tmp_i_cast_fu_777_p1 = $signed(tmp_39_i_fu_767_p4);
  assign tmp_i_fu_581_p2 = $signed(reg_481) * $signed(reg_477);
  assign tmp_s_fu_566_p1 = tmp_1_cast_fu_557_p4;
  assign wd1_2_fu_1364_p4 = { { nbl_assign_6_fu_1346_p3[10:6] } };
  assign wd1_fu_742_p4 = { { nbl_assign_5_fu_724_p3[10:6] } };
  assign wd2_15_cast_fu_983_p1 = $signed(tmp_55_fu_975_p3);
  assign wd2_16_cast_fu_1096_p1 = $signed(tmp_21_i_reg_2020);
  assign wd2_21_cast_fu_1551_p1 = $signed(tmp_58_fu_1543_p3);
  assign wd2_22_cast_fu_1680_p1 = $signed(tmp_21_i2_reg_2149);
  assign wd2_4_fu_949_p2 = 32'd0 - wd2_fu_936_p2;
  assign wd2_5_fu_1504_p2 = dec_ah1_i << 32'd2;
  assign wd2_6_fu_1517_p2 = 32'd0 - wd2_5_fu_1504_p2;
  assign wd2_fu_936_p2 = dec_al1_i << 32'd2;
  assign wd3_0_apl1_i2_fu_1747_p3 = (tmp_6_i2_fu_1742_p2[0:0] === 1'b1)? apl1_18_cast_fu_1738_p1 : apl1_13_reg_2170;
  assign wd3_0_apl1_i_fu_1145_p3 = (tmp_6_i_fu_1140_p2[0:0] === 1'b1)? apl1_17_cast_fu_1136_p1 : apl1_reg_2031;
  assign wd3_5_fu_1424_p2 = ilb_table_q0 >> tmp_9_i5_cast_cast_fu_1420_p1;
  assign wd3_fu_834_p2 = ilb_table_q0 >> tmp_9_i_cast_cast_fu_830_p1;
  assign wd_cast_fu_618_p1 = tmp_32_i_fu_608_p4;
  assign wd_fu_1256_p1 = tmp_36_i_fu_1246_p4;
  assign wl_code_table_address0 = tmp_s_fu_566_p1;
  assign wl_code_table_load_c_fu_622_p0 = wl_code_table_q0;
  assign wl_code_table_load_c_fu_622_p1 = wl_code_table_load_c_fu_622_p0;
  assign xd_fu_1819_p2 = $signed(rl_cast_reg_2057) - $signed(rh_fu_1801_p2);
  assign xs_fu_1824_p2 = $signed(rh_fu_1801_p2) + $signed(rl_cast_reg_2057);
  assign zl_5_fu_587_p2 = tmp_i_reg_1928 + zl1_i_reg_378;
  assign zl_6_fu_1302_p2 = tmp_i8_33_reg_2096 + zl1_i2_reg_399;
  assign zl_fu_499_p2 = $signed(reg_477) * $signed(reg_481);
  assign temp140 = temp142 * temp143;
  assign temp143 = (working_key[39] == 1'b1)? dec_nbl_i + dec_detl_i : dec_al2_i + dec_del_dltx_q0;
  assign temp142 = (working_key[40] == 1'b1)? dec_al2_i + dec_rlt2_i : dec_del_dhx_q1 + ih_i;
  assign temp144 = temp146 * temp147;
  assign temp147 = (working_key[42] == 1'b1)? dec_detl_i + dec_deth_i : ih_i + dec_del_bph_q0;
  assign temp146 = (working_key[43] == 1'b1)? dec_del_dhx_q1 + dec_plt1_i : accumc_q0 + ih_i;
  assign temp148 = temp150 * temp151;
  assign temp151 = (working_key[45] == 1'b1)? dec_del_bpl_q0 + dec_nbh_i : dec_nbl_i + dec_ph1_i;
  assign temp150 = (working_key[46] == 1'b1)? dec_plt2_i + accumc_q0 : dec_ah2_i + ih_i;
  assign temp152 = temp154 * temp155;
  assign temp155 = (working_key[48] == 1'b1)? dec_del_bpl_q0 + dec_detl_i : dec_al2_i + accumc_q0;
  assign temp154 = (working_key[49] == 1'b1)? dec_nbh_i + dec_deth_i : dec_nbh_i + dec_detl_i;
  assign temp156 = temp158 * temp159;
  assign temp159 = (working_key[51] == 1'b1)? dec_del_dltx_q0 + dec_del_bpl_q0 : dec_del_dltx_q1 + dec_plt2_i;
  assign temp158 = (working_key[52] == 1'b1)? dec_del_dhx_q1 + dec_deth_i : dec_al2_i + dec_al1_i;
  assign temp160 = temp162 * temp163;
  assign temp163 = (working_key[54] == 1'b1)? il + dec_al2_i : dec_rh2_i + dec_nbh_i;
  assign temp162 = (working_key[55] == 1'b1)? dec_al2_i + dec_ah2_i : accumd_q0 + dec_del_dhx_q0;
  assign temp164 = temp166 * temp167;
  assign temp167 = (working_key[57] == 1'b1)? input_r + dec_del_bph_q0 : dec_ah1_i + input_r;
  assign temp166 = (working_key[58] == 1'b1)? dec_del_dhx_q1 + dec_deth_i : dec_ah1_i + dec_del_dltx_q1;
  assign temp168 = temp170 * temp171;
  assign temp171 = (working_key[59] == 1'b1)? dec_ph1_i + dec_detl_i : dec_al2_i + dec_del_bpl_q0;
  assign temp170 = (working_key[60] == 1'b1)? dec_nbh_i + dec_detl_i : dec_rlt2_i + accumc_q0;
  assign temp172 = temp174 * temp175;
  assign temp175 = (working_key[61] == 1'b1)? dec_deth_i + ih_i : dec_del_dhx_q0 + accumd_q0;
  assign temp174 = (working_key[62] == 1'b1)? dec_ph1_i + dec_nbl_i : input_r + dec_del_dltx_q1;
  assign temp176 = temp178 * temp179;
  assign temp179 = (working_key[63] == 1'b1)? dec_ah2_i + dec_del_bph_q0 : dec_plt1_i + dec_ah1_i;
  assign temp178 = (working_key[64] == 1'b1)? dec_plt1_i + dec_ah1_i : dec_rlt2_i + dec_del_dhx_q1;

endmodule


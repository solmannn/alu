
module decode_0_obf
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  input_r,
  ih_i,
  ih_o,
  ih_o_ap_vld,
  dec_del_bpl_address0,
  dec_del_bpl_ce0,
  dec_del_bpl_we0,
  dec_del_bpl_d0,
  dec_del_bpl_q0,
  dec_del_dltx_address0,
  dec_del_dltx_ce0,
  dec_del_dltx_we0,
  dec_del_dltx_d0,
  dec_del_dltx_q0,
  dec_del_dltx_address1,
  dec_del_dltx_ce1,
  dec_del_dltx_we1,
  dec_del_dltx_d1,
  dec_del_dltx_q1,
  dec_rlt1_i,
  dec_rlt1_o,
  dec_rlt1_o_ap_vld,
  dec_al1_i,
  dec_al1_o,
  dec_al1_o_ap_vld,
  dec_rlt2_i,
  dec_rlt2_o,
  dec_rlt2_o_ap_vld,
  dec_al2_i,
  dec_al2_o,
  dec_al2_o_ap_vld,
  dec_detl_i,
  dec_detl_o,
  dec_detl_o_ap_vld,
  il,
  dec_nbl_i,
  dec_nbl_o,
  dec_nbl_o_ap_vld,
  dec_plt1_i,
  dec_plt1_o,
  dec_plt1_o_ap_vld,
  dec_plt2_i,
  dec_plt2_o,
  dec_plt2_o_ap_vld,
  dec_del_bph_address0,
  dec_del_bph_ce0,
  dec_del_bph_we0,
  dec_del_bph_d0,
  dec_del_bph_q0,
  dec_del_dhx_address0,
  dec_del_dhx_ce0,
  dec_del_dhx_we0,
  dec_del_dhx_d0,
  dec_del_dhx_q0,
  dec_del_dhx_address1,
  dec_del_dhx_ce1,
  dec_del_dhx_we1,
  dec_del_dhx_d1,
  dec_del_dhx_q1,
  dec_rh1_i,
  dec_rh1_o,
  dec_rh1_o_ap_vld,
  dec_ah1_i,
  dec_ah1_o,
  dec_ah1_o_ap_vld,
  dec_rh2_i,
  dec_rh2_o,
  dec_rh2_o_ap_vld,
  dec_ah2_i,
  dec_ah2_o,
  dec_ah2_o_ap_vld,
  dec_deth_i,
  dec_deth_o,
  dec_deth_o_ap_vld,
  dec_nbh_i,
  dec_nbh_o,
  dec_nbh_o_ap_vld,
  dec_ph1_i,
  dec_ph1_o,
  dec_ph1_o_ap_vld,
  dec_ph2_i,
  dec_ph2_o,
  dec_ph2_o_ap_vld,
  accumc_address0,
  accumc_ce0,
  accumc_we0,
  accumc_d0,
  accumc_q0,
  accumd_address0,
  accumd_ce0,
  accumd_we0,
  accumd_d0,
  accumd_q0,
  locking_key
);

  parameter ap_ST_fsm_state1 = 29'd1;
  parameter ap_ST_fsm_state2 = 29'd2;
  parameter ap_ST_fsm_state3 = 29'd4;
  parameter ap_ST_fsm_state4 = 29'd8;
  parameter ap_ST_fsm_state5 = 29'd16;
  parameter ap_ST_fsm_state6 = 29'd32;
  parameter ap_ST_fsm_state7 = 29'd64;
  parameter ap_ST_fsm_state8 = 29'd128;
  parameter ap_ST_fsm_state9 = 29'd256;
  parameter ap_ST_fsm_state10 = 29'd512;
  parameter ap_ST_fsm_state11 = 29'd1024;
  parameter ap_ST_fsm_state12 = 29'd2048;
  parameter ap_ST_fsm_state13 = 29'd4096;
  parameter ap_ST_fsm_state14 = 29'd8192;
  parameter ap_ST_fsm_state15 = 29'd16384;
  parameter ap_ST_fsm_state16 = 29'd32768;
  parameter ap_ST_fsm_state17 = 29'd65536;
  parameter ap_ST_fsm_state18 = 29'd131072;
  parameter ap_ST_fsm_state19 = 29'd262144;
  parameter ap_ST_fsm_state20 = 29'd524288;
  parameter ap_ST_fsm_state21 = 29'd1048576;
  parameter ap_ST_fsm_state22 = 29'd2097152;
  parameter ap_ST_fsm_state23 = 29'd4194304;
  parameter ap_ST_fsm_state24 = 29'd8388608;
  parameter ap_ST_fsm_state25 = 29'd16777216;
  parameter ap_ST_fsm_state26 = 29'd33554432;
  parameter ap_ST_fsm_state27 = 29'd67108864;
  parameter ap_ST_fsm_state28 = 29'd134217728;
  parameter ap_ST_fsm_state29 = 29'd268435456;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  input [31:0] input_r;
  input [31:0] ih_i;
  output [31:0] ih_o;
  output ih_o_ap_vld;
  output [2:0] dec_del_bpl_address0;
  output dec_del_bpl_ce0;
  output dec_del_bpl_we0;
  output [31:0] dec_del_bpl_d0;
  input [31:0] dec_del_bpl_q0;
  output [2:0] dec_del_dltx_address0;
  output dec_del_dltx_ce0;
  output dec_del_dltx_we0;
  output [31:0] dec_del_dltx_d0;
  input [31:0] dec_del_dltx_q0;
  output [2:0] dec_del_dltx_address1;
  output dec_del_dltx_ce1;
  output dec_del_dltx_we1;
  output [31:0] dec_del_dltx_d1;
  input [31:0] dec_del_dltx_q1;
  input [31:0] dec_rlt1_i;
  output [31:0] dec_rlt1_o;
  output dec_rlt1_o_ap_vld;
  input [31:0] dec_al1_i;
  output [31:0] dec_al1_o;
  output dec_al1_o_ap_vld;
  input [31:0] dec_rlt2_i;
  output [31:0] dec_rlt2_o;
  output dec_rlt2_o_ap_vld;
  input [31:0] dec_al2_i;
  output [31:0] dec_al2_o;
  output dec_al2_o_ap_vld;
  input [14:0] dec_detl_i;
  output [14:0] dec_detl_o;
  output dec_detl_o_ap_vld;
  input [5:0] il;
  input [31:0] dec_nbl_i;
  output [31:0] dec_nbl_o;
  output dec_nbl_o_ap_vld;
  input [31:0] dec_plt1_i;
  output [31:0] dec_plt1_o;
  output dec_plt1_o_ap_vld;
  input [31:0] dec_plt2_i;
  output [31:0] dec_plt2_o;
  output dec_plt2_o_ap_vld;
  output [2:0] dec_del_bph_address0;
  output dec_del_bph_ce0;
  output dec_del_bph_we0;
  output [31:0] dec_del_bph_d0;
  input [31:0] dec_del_bph_q0;
  output [2:0] dec_del_dhx_address0;
  output dec_del_dhx_ce0;
  output dec_del_dhx_we0;
  output [31:0] dec_del_dhx_d0;
  input [31:0] dec_del_dhx_q0;
  output [2:0] dec_del_dhx_address1;
  output dec_del_dhx_ce1;
  output dec_del_dhx_we1;
  output [31:0] dec_del_dhx_d1;
  input [31:0] dec_del_dhx_q1;
  input [31:0] dec_rh1_i;
  output [31:0] dec_rh1_o;
  output dec_rh1_o_ap_vld;
  input [31:0] dec_ah1_i;
  output [31:0] dec_ah1_o;
  output dec_ah1_o_ap_vld;
  input [31:0] dec_rh2_i;
  output [31:0] dec_rh2_o;
  output dec_rh2_o_ap_vld;
  input [31:0] dec_ah2_i;
  output [31:0] dec_ah2_o;
  output dec_ah2_o_ap_vld;
  input [14:0] dec_deth_i;
  output [14:0] dec_deth_o;
  output dec_deth_o_ap_vld;
  input [31:0] dec_nbh_i;
  output [31:0] dec_nbh_o;
  output dec_nbh_o_ap_vld;
  input [31:0] dec_ph1_i;
  output [31:0] dec_ph1_o;
  output dec_ph1_o_ap_vld;
  input [31:0] dec_ph2_i;
  output [31:0] dec_ph2_o;
  output dec_ph2_o_ap_vld;
  output [3:0] accumc_address0;
  output accumc_ce0;
  output accumc_we0;
  output [31:0] accumc_d0;
  input [31:0] accumc_q0;
  output [3:0] accumd_address0;
  output accumd_ce0;
  output accumd_we0;
  output [31:0] accumd_d0;
  input [31:0] accumd_q0;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [31:0] ih_o;
  reg ih_o_ap_vld;
  reg [2:0] dec_del_bpl_address0;
  reg dec_del_bpl_ce0;
  reg dec_del_bpl_we0;
  reg [2:0] dec_del_dltx_address0;
  reg dec_del_dltx_ce0;
  reg dec_del_dltx_we0;
  reg dec_del_dltx_ce1;
  reg dec_del_dltx_we1;
  reg [31:0] dec_rlt1_o;
  reg dec_rlt1_o_ap_vld;
  reg [31:0] dec_al1_o;
  reg dec_al1_o_ap_vld;
  reg [31:0] dec_rlt2_o;
  reg dec_rlt2_o_ap_vld;
  reg [31:0] dec_al2_o;
  reg dec_al2_o_ap_vld;
  reg [14:0] dec_detl_o;
  reg dec_detl_o_ap_vld;
  reg [31:0] dec_nbl_o;
  reg dec_nbl_o_ap_vld;
  reg [31:0] dec_plt1_o;
  reg dec_plt1_o_ap_vld;
  reg [31:0] dec_plt2_o;
  reg dec_plt2_o_ap_vld;
  reg [2:0] dec_del_bph_address0;
  reg dec_del_bph_ce0;
  reg dec_del_bph_we0;
  reg [2:0] dec_del_dhx_address0;
  reg dec_del_dhx_ce0;
  reg dec_del_dhx_we0;
  reg dec_del_dhx_ce1;
  reg dec_del_dhx_we1;
  reg [31:0] dec_rh1_o;
  reg dec_rh1_o_ap_vld;
  reg [31:0] dec_ah1_o;
  reg dec_ah1_o_ap_vld;
  reg [31:0] dec_rh2_o;
  reg dec_rh2_o_ap_vld;
  reg [31:0] dec_ah2_o;
  reg dec_ah2_o_ap_vld;
  reg [14:0] dec_deth_o;
  reg dec_deth_o_ap_vld;
  reg [31:0] dec_nbh_o;
  reg dec_nbh_o_ap_vld;
  reg [31:0] dec_ph1_o;
  reg dec_ph1_o_ap_vld;
  reg [31:0] dec_ph2_o;
  reg dec_ph2_o_ap_vld;
  reg [3:0] accumc_address0;
  reg accumc_ce0;
  reg accumc_we0;
  reg [31:0] accumc_d0;
  reg [3:0] accumd_address0;
  reg accumd_ce0;
  reg accumd_we0;
  reg [31:0] accumd_d0;
  reg [28:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  wire [3:0] qq4_code4_table_address0;
  reg qq4_code4_table_ce0;
  wire [15:0] qq4_code4_table_q0;
  reg [31:0] dec_dlt;
  wire [5:0] qq6_code6_table_address0;
  reg qq6_code6_table_ce0;
  wire [15:0] qq6_code6_table_q0;
  wire [3:0] wl_code_table_address0;
  reg wl_code_table_ce0;
  wire [12:0] wl_code_table_q0;
  reg [4:0] ilb_table_address0;
  reg ilb_table_ce0;
  wire [11:0] ilb_table_q0;
  reg [31:0] dec_plt;
  reg [31:0] dec_dh;
  reg [31:0] dec_ph;
  reg signed [31:0] reg_477;
  wire ap_CS_fsm_state2;
  wire ap_CS_fsm_state6;
  reg signed [31:0] reg_481;
  reg signed [31:0] reg_485;
  wire ap_CS_fsm_state14;
  wire ap_CS_fsm_state18;
  reg signed [31:0] reg_489;
  wire [31:0] zl_fu_499_p2;
  reg [31:0] zl_reg_1885;
  wire ap_CS_fsm_state3;
  wire ap_CS_fsm_state4;
  wire [2:0] p_01_rec_i_fu_539_p2;
  reg [2:0] p_01_rec_i_reg_1895;
  wire ap_CS_fsm_state5;
  wire [0:0] exitcond3_fu_551_p2;
  wire [31:0] tmp_i_fu_581_p2;
  reg [31:0] tmp_i_reg_1928;
  wire ap_CS_fsm_state7;
  wire [31:0] zl_5_fu_587_p2;
  wire ap_CS_fsm_state8;
  reg signed [15:0] qq4_code4_table_load_reg_1938;
  wire ap_CS_fsm_state9;
  reg signed [15:0] qq6_code6_table_load_reg_1943;
  wire [24:0] nbl_assign_4_cast_fu_636_p2;
  reg [24:0] nbl_assign_4_cast_reg_1948;
  reg [0:0] tmp_73_reg_1953;
  wire [31:0] pl_fu_654_p2;
  reg [31:0] pl_reg_1958;
  wire ap_CS_fsm_state10;
  wire [31:0] tmp_i1_fu_660_p2;
  reg [31:0] tmp_i1_reg_1963;
  wire signed [15:0] tmp_70_fu_677_p4;
  reg signed [15:0] tmp_70_reg_1968;
  reg [15:0] tmp_71_reg_1974;
  reg [3:0] wd2_cast_reg_1979;
  wire signed [16:0] tmp_43_fu_809_p1;
  reg signed [16:0] tmp_43_reg_1989;
  wire ap_CS_fsm_state11;
  wire [18:0] rl_fu_819_p2;
  reg [18:0] rl_reg_1994;
  wire [31:0] tmp_i8_fu_904_p2;
  reg [31:0] tmp_i8_reg_1999;
  wire ap_CS_fsm_state12;
  wire grp_upzero_fu_442_ap_ready;
  wire grp_upzero_fu_442_ap_done;
  wire [31:0] tmp_5_i_fu_910_p2;
  reg [31:0] tmp_5_i_reg_2004;
  reg [0:0] tmp_81_reg_2009;
  wire [26:0] apl2_fu_1038_p2;
  reg [26:0] apl2_reg_2014;
  wire ap_CS_fsm_state13;
  reg [23:0] tmp_21_i_reg_2020;
  wire signed [14:0] apl2_assign_fu_1088_p3;
  reg signed [14:0] apl2_assign_reg_2025;
  wire [24:0] apl1_fu_1112_p2;
  reg [24:0] apl1_reg_2031;
  wire [15:0] tmp_82_fu_1152_p1;
  reg [15:0] tmp_82_reg_2037;
  wire ap_CS_fsm_state15;
  wire signed [15:0] apl1_11_fu_1156_p2;
  reg signed [15:0] apl1_11_reg_2042;
  wire [0:0] tmp_7_i_fu_1166_p2;
  reg [0:0] tmp_7_i_reg_2047;
  wire [31:0] grp_fu_493_p2;
  reg [31:0] zl_4_reg_2052;
  wire signed [31:0] rl_cast_fu_1172_p1;
  reg signed [31:0] rl_cast_reg_2057;
  wire ap_CS_fsm_state16;
  wire [2:0] p_01_rec_i2_fu_1190_p2;
  reg [2:0] p_01_rec_i2_reg_2063;
  wire ap_CS_fsm_state17;
  wire signed [31:0] tmp_14_fu_1216_p6;
  reg signed [31:0] tmp_14_reg_2081;
  wire [0:0] exitcond2_fu_1202_p2;
  wire [30:0] nbh_assign_2_cast_fu_1288_p2;
  reg [30:0] nbh_assign_2_cast_reg_2086;
  reg [0:0] tmp_86_reg_2091;
  reg [31:0] tmp_i8_33_reg_2096;
  wire ap_CS_fsm_state19;
  wire [31:0] zl_6_fu_1302_p2;
  wire ap_CS_fsm_state20;
  reg signed [16:0] tmp_50_reg_2106;
  wire ap_CS_fsm_state21;
  reg [3:0] wd2_17_cast_reg_2113;
  wire signed [18:0] tmp_i19_cast_fu_1399_p1;
  reg signed [18:0] tmp_i19_cast_reg_2123;
  wire ap_CS_fsm_state22;
  wire [31:0] tmp_i3_fu_1472_p2;
  reg [31:0] tmp_i3_reg_2128;
  wire ap_CS_fsm_state23;
  wire [31:0] tmp_5_i5_fu_1478_p2;
  reg [31:0] tmp_5_i5_reg_2133;
  reg [0:0] tmp_94_reg_2138;
  wire [26:0] apl2_2_fu_1606_p2;
  reg [26:0] apl2_2_reg_2143;
  wire ap_CS_fsm_state24;
  reg [23:0] tmp_21_i2_reg_2149;
  wire [31:0] pl_2_fu_1638_p2;
  reg [31:0] pl_2_reg_2154;
  wire ap_CS_fsm_state25;
  wire [31:0] tmp_i4_fu_1644_p2;
  reg [31:0] tmp_i4_reg_2159;
  wire signed [14:0] apl2_assign_2_fu_1672_p3;
  reg signed [14:0] apl2_assign_2_reg_2164;
  wire [24:0] apl1_13_fu_1696_p2;
  reg [24:0] apl1_13_reg_2170;
  wire [15:0] tmp_95_fu_1754_p1;
  reg [15:0] tmp_95_reg_2176;
  wire ap_CS_fsm_state26;
  wire signed [15:0] apl1_15_fu_1758_p2;
  reg signed [15:0] apl1_15_reg_2181;
  wire [0:0] tmp_7_i2_fu_1768_p2;
  reg [0:0] tmp_7_i2_reg_2186;
  wire [18:0] tmp8_fu_1774_p2;
  reg [18:0] tmp8_reg_2191;
  wire [31:0] xd_fu_1819_p2;
  reg [31:0] xd_reg_2196;
  wire ap_CS_fsm_state27;
  wire [31:0] xs_fu_1824_p2;
  reg [31:0] xs_reg_2201;
  reg [3:0] accumc_addr_reg_2206;
  wire ap_CS_fsm_state28;
  reg [3:0] accumd_addr_reg_2211;
  wire [4:0] p_rec_fu_1841_p2;
  reg [4:0] p_rec_reg_2216;
  wire [3:0] i_fu_1865_p2;
  reg [3:0] i_reg_2234;
  wire grp_upzero_fu_442_ap_start;
  wire grp_upzero_fu_442_ap_idle;
  reg [16:0] grp_upzero_fu_442_dlt;
  wire [2:0] grp_upzero_fu_442_dlti_address0;
  wire grp_upzero_fu_442_dlti_ce0;
  wire grp_upzero_fu_442_dlti_we0;
  wire [31:0] grp_upzero_fu_442_dlti_d0;
  reg [31:0] grp_upzero_fu_442_dlti_q0;
  wire [2:0] grp_upzero_fu_442_dlti_address1;
  wire grp_upzero_fu_442_dlti_ce1;
  wire grp_upzero_fu_442_dlti_we1;
  wire [31:0] grp_upzero_fu_442_dlti_d1;
  reg [31:0] grp_upzero_fu_442_dlti_q1;
  wire [2:0] grp_upzero_fu_442_bli_address0;
  wire grp_upzero_fu_442_bli_ce0;
  wire grp_upzero_fu_442_bli_we0;
  wire [31:0] grp_upzero_fu_442_bli_d0;
  reg [31:0] grp_upzero_fu_442_bli_q0;
  reg [31:0] zl1_i_reg_378;
  reg [2:0] dlt_pn_rec_i_reg_388;
  reg [31:0] zl1_i2_reg_399;
  reg [2:0] dlt_pn_rec_i2_reg_409;
  reg [4:0] ad_ptr_1_rec_reg_420;
  wire ap_CS_fsm_state29;
  reg [3:0] i_1_reg_431;
  reg grp_upzero_fu_442_ap_start_reg;
  wire [63:0] p_01_rec_i_cast_fu_545_p1;
  wire [63:0] tmp_s_fu_566_p1;
  wire [63:0] tmp_45_fu_576_p1;
  wire [63:0] tmp_i2_fu_762_p1;
  wire [63:0] p_01_rec_i2_cast_fu_1196_p1;
  wire [63:0] tmp_i6_fu_1384_p1;
  wire [63:0] ac_ptr_0_sum_cast_fu_1835_p1;
  wire [63:0] ad_ptr_0_sum7_cast_fu_1853_p1;
  wire signed [31:0] tmp_44_fu_686_p1;
  wire signed [31:0] tmp_64_cast_fu_860_p1;
  wire signed [31:0] tmp_51_fu_1403_p1;
  wire signed [31:0] tmp_70_cast_fu_1450_p1;
  wire signed [31:0] ih_assign_fu_529_p1;
  wire [31:0] nbl_assign_5_cast_fu_732_p1;
  wire [14:0] tmp_10_i_fu_840_p3;
  wire [31:0] dec_rlt_fu_874_p2;
  wire signed [31:0] apl2_assign_cast_fu_1118_p1;
  wire signed [31:0] apl1_12_cast_fu_1180_p1;
  wire [31:0] nbl_assign_6_cast_fu_1354_p1;
  wire [14:0] tmp_10_i2_fu_1430_p3;
  wire signed [31:0] apl2_assign_2_cast_fu_1720_p1;
  wire signed [31:0] apl1_16_cast_fu_1784_p1;
  wire [31:0] rh_fu_1801_p2;
  wire [0:0] exitcond_fu_1859_p2;
  wire [25:0] tmp_41_fu_519_p4;
  wire [3:0] tmp_1_cast_fu_557_p4;
  wire [31:0] tmp_72_fu_596_p2;
  wire [31:0] tmp_i7_fu_602_p2;
  wire signed [24:0] tmp_32_i_fu_608_p4;
  wire signed [12:0] wl_code_table_load_c_fu_622_p0;
  wire signed [12:0] tmp_13_fu_626_p0;
  wire signed [25:0] wd_cast_fu_618_p1;
  wire signed [25:0] wl_code_table_load_c_fu_622_p1;
  wire signed [24:0] tmp_13_fu_626_p1;
  wire [25:0] nbl_assign_4_fu_630_p2;
  wire signed [31:0] pl_fu_654_p0;
  wire signed [31:0] pl_fu_654_p1;
  wire signed [31:0] tmp_i1_fu_660_p0;
  wire signed [31:0] tmp_i1_fu_660_p1;
  wire signed [30:0] tmp_42_fu_1871_p2;
  wire signed [30:0] tmp_46_fu_1878_p2;
  wire [24:0] p_i_fu_708_p3;
  wire [0:0] tmp_18_i_fu_718_p2;
  wire [14:0] tmp_74_fu_714_p1;
  wire [14:0] nbl_assign_5_fu_724_p3;
  wire [4:0] wd1_fu_742_p4;
  wire [17:0] tmp_39_i_fu_767_p4;
  wire [31:0] tmp_i_31_fu_781_p2;
  wire [16:0] tmp_41_i_fu_785_p4;
  wire signed [18:0] tmp_20_i_cast_fu_795_p1;
  wire signed [18:0] tmp_i_cast_fu_777_p1;
  wire signed [18:0] dec_sl_fu_799_p2;
  wire signed [18:0] dl_cast_fu_816_p1;
  wire [3:0] tmp_9_i_fu_825_p2;
  wire [11:0] tmp_9_i_cast_cast_fu_830_p1;
  wire [11:0] wd3_fu_834_p2;
  wire signed [18:0] tmp_59_cast_fu_813_p1;
  wire [18:0] tmp_48_fu_854_p2;
  wire signed [31:0] dec_sl_cast_fu_805_p1;
  wire signed [31:0] tmp_i8_fu_904_p0;
  wire signed [31:0] tmp_i8_fu_904_p1;
  wire signed [31:0] tmp_5_i_fu_910_p0;
  wire signed [31:0] tmp_5_i_fu_910_p1;
  wire [31:0] wd2_fu_936_p2;
  wire [31:0] wd2_4_fu_949_p2;
  wire [0:0] tmp_76_fu_942_p3;
  wire [24:0] tmp_54_fu_965_p4;
  wire [24:0] tmp_53_fu_955_p4;
  wire [24:0] tmp_55_fu_975_p3;
  wire [0:0] tmp_77_fu_987_p3;
  wire [31:0] tmp_78_fu_1002_p2;
  wire [31:0] tmp_9_i4_fu_1008_p2;
  wire [24:0] tmp_19_i_fu_1014_p4;
  wire signed [25:0] wd2_15_cast_fu_983_p1;
  wire signed [25:0] tmp_1_i_cast_fu_1024_p1;
  wire [25:0] tmp4_fu_1028_p2;
  wire [26:0] tmp_8_i_cast_cast_fu_994_p3;
  wire signed [26:0] tmp4_cast_fu_1034_p1;
  wire [31:0] tmp_80_fu_1044_p2;
  wire [31:0] tmp_i9_fu_1050_p2;
  wire [0:0] tmp_2_i_fu_1066_p2;
  wire [26:0] p_i4_fu_1071_p3;
  wire [0:0] tmp_3_i_fu_1082_p2;
  wire [14:0] tmp_79_fu_1078_p1;
  wire signed [24:0] wd2_16_cast_fu_1096_p1;
  wire [24:0] tmp_4_i_cast_cast_fu_1099_p3;
  wire [24:0] tmp5_fu_1106_p2;
  wire [14:0] apl1_17_fu_1127_p2;
  wire [24:0] apl1_17_cast_fu_1136_p1;
  wire [0:0] tmp_6_i_fu_1140_p2;
  wire [24:0] wd3_0_apl1_i_fu_1145_p3;
  wire [15:0] apl1_17_cast1_fu_1132_p1;
  wire signed [24:0] apl1_11_cast_fu_1162_p1;
  wire [15:0] apl1_12_fu_1175_p3;
  wire [1:0] tmp_83_fu_1212_p1;
  wire [31:0] tmp_84_fu_1234_p2;
  wire [31:0] tmp_i2_35_fu_1240_p2;
  wire signed [24:0] tmp_36_i_fu_1246_p4;
  wire [31:0] tmp_15_fu_1260_p6;
  wire signed [31:0] wd_fu_1256_p1;
  wire signed [30:0] tmp_16_fu_1274_p1;
  wire [30:0] tmp_85_fu_1278_p1;
  wire [31:0] nbh_assign_2_fu_1282_p2;
  wire [14:0] tmp_49_fu_1315_p0;
  wire [31:0] tmp_49_fu_1315_p2;
  wire [30:0] p_i5_fu_1330_p3;
  wire [0:0] tmp_19_i3_fu_1340_p2;
  wire [14:0] tmp_87_fu_1336_p1;
  wire [14:0] nbl_assign_6_fu_1346_p3;
  wire [4:0] wd1_2_fu_1364_p4;
  wire [17:0] tmp_39_i2_fu_1389_p4;
  wire [3:0] tmp_9_i5_fu_1415_p2;
  wire [11:0] tmp_9_i5_cast_cast_fu_1420_p1;
  wire [11:0] wd3_5_fu_1424_p2;
  wire signed [18:0] tmp_69_cast_fu_1406_p1;
  wire [18:0] tmp_52_fu_1444_p2;
  wire signed [31:0] tmp_i3_fu_1472_p0;
  wire signed [31:0] tmp_i3_fu_1472_p1;
  wire signed [31:0] tmp_5_i5_fu_1478_p0;
  wire signed [31:0] tmp_5_i5_fu_1478_p1;
  wire [31:0] wd2_5_fu_1504_p2;
  wire [31:0] wd2_6_fu_1517_p2;
  wire [0:0] tmp_89_fu_1510_p3;
  wire [24:0] tmp_57_fu_1533_p4;
  wire [24:0] tmp_56_fu_1523_p4;
  wire [24:0] tmp_58_fu_1543_p3;
  wire [0:0] tmp_90_fu_1555_p3;
  wire [31:0] tmp_91_fu_1570_p2;
  wire [31:0] tmp_9_i6_fu_1576_p2;
  wire [24:0] tmp_19_i4_fu_1582_p4;
  wire signed [25:0] tmp_1_i2_cast_fu_1592_p1;
  wire signed [25:0] wd2_21_cast_fu_1551_p1;
  wire [25:0] tmp6_fu_1596_p2;
  wire signed [26:0] tmp6_cast_fu_1602_p1;
  wire [26:0] tmp_8_i2_cast_cast_fu_1562_p3;
  wire [31:0] tmp_93_fu_1612_p2;
  wire [31:0] tmp_i4_36_fu_1618_p2;
  wire signed [31:0] pl_2_fu_1638_p0;
  wire signed [31:0] pl_2_fu_1638_p1;
  wire signed [31:0] tmp_i4_fu_1644_p0;
  wire signed [31:0] tmp_i4_fu_1644_p1;
  wire [0:0] tmp_2_i2_fu_1650_p2;
  wire [26:0] p_i6_fu_1655_p3;
  wire [0:0] tmp_3_i2_fu_1666_p2;
  wire [14:0] tmp_92_fu_1662_p1;
  wire signed [24:0] wd2_22_cast_fu_1680_p1;
  wire [24:0] tmp7_fu_1690_p2;
  wire [24:0] tmp_4_i2_cast_cast_fu_1683_p3;
  wire [31:0] tmp_i1_34_fu_1702_p2;
  wire [16:0] tmp_41_i2_fu_1706_p4;
  wire [14:0] apl1_18_fu_1729_p2;
  wire [24:0] apl1_18_cast_fu_1738_p1;
  wire [0:0] tmp_6_i2_fu_1742_p2;
  wire [24:0] wd3_0_apl1_i2_fu_1747_p3;
  wire [15:0] apl1_18_cast9_fu_1734_p1;
  wire signed [24:0] apl1_15_cast_fu_1764_p1;
  wire signed [18:0] tmp_20_i5_cast_fu_1716_p1;
  wire [15:0] apl1_16_fu_1779_p3;
  wire signed [31:0] tmp8_cast_fu_1798_p1;
  wire [4:0] ac_ptr_0_sum_fu_1829_p2;
  wire [4:0] ad_ptr_0_sum7_fu_1847_p2;
  wire [14:0] tmp_42_fu_1871_p1;
  wire [30:0] extLd_cast_fu_670_p1;
  wire [14:0] tmp_46_fu_1878_p1;
  reg [28:0] ap_NS_fsm;
  wire [31:0] tmp_49_fu_1315_p00;
  wire [31:0] Const_197;
  wire [31:0] Const_198;
  wire [31:0] Const_199;
  wire [31:0] Const_200;
  wire [31:0] Const_201;
  wire [31:0] Const_202;
  wire [31:0] Const_203;
  wire [31:0] Const_204;
  wire Const_205;
  wire [4:0] Const_206;
  wire Const_207;
  wire Const_208;
  wire Const_209;
  wire [2:0] Const_210;
  wire Const_211;
  wire Const_212;
  wire [2:0] Const_213;
  wire Const_214;
  wire [3:0] Const_215;
  wire Const_216;
  wire Const_217;
  wire Const_218;
  wire Const_219;
  wire Const_220;
  wire Const_221;
  wire Const_222;
  wire Const_223;
  wire Const_224;
  wire Const_225;
  wire Const_226;
  wire Const_227;
  wire Const_228;
  wire Const_229;
  wire Const_230;
  wire Const_231;
  wire Const_232;
  wire Const_233;
  wire Const_234;
  wire Const_235;
  wire Const_236;
  wire Const_237;
  wire Const_238;
  wire Const_239;
  wire Const_240;
  wire Const_241;
  wire Const_242;
  wire Const_243;
  wire Const_244;
  wire Const_245;
  wire Const_246;
  wire Const_247;
  wire Const_248;
  wire Const_249;
  wire Const_250;
  wire Const_251;
  wire Const_252;
  wire [3:0] Const_253;
  wire Const_254;
  wire Const_255;
  wire Const_256;
  wire Const_257;
  wire Const_258;
  wire Const_259;
  wire Const_260;
  wire Const_261;
  wire Const_262;
  wire Const_263;
  wire Const_264;
  wire Const_265;
  wire Const_266;
  wire Const_267;
  wire Const_268;
  wire Const_269;
  wire Const_270;
  wire Const_271;
  wire Const_272;
  wire Const_273;
  wire [3:0] Const_274;
  wire Const_275;
  wire Const_276;
  wire Const_277;
  wire Const_278;
  wire Const_279;
  wire Const_280;
  wire Const_281;
  wire Const_282;
  wire Const_283;
  wire Const_284;
  wire Const_285;
  wire Const_286;
  wire Const_287;
  wire Const_288;
  wire Const_289;
  wire Const_290;
  wire Const_291;
  wire Const_292;
  wire Const_293;
  wire Const_294;
  wire Const_295;
  wire Const_296;
  wire Const_297;
  wire Const_298;
  wire Const_299;
  wire Const_300;
  wire Const_301;
  wire Const_302;
  wire Const_303;
  wire Const_304;
  wire Const_305;
  wire Const_306;
  wire Const_307;
  wire Const_308;
  wire Const_309;
  wire Const_310;
  wire Const_311;
  wire Const_312;
  wire Const_313;
  wire Const_314;
  wire Const_315;
  wire Const_316;
  wire Const_317;
  wire Const_318;
  wire Const_319;
  wire Const_320;
  wire Const_321;
  wire Const_322;
  wire Const_323;
  wire [2:0] Const_324;
  wire Const_325;
  wire Const_326;
  wire Const_327;
  wire Const_328;
  wire Const_329;
  wire Const_330;
  wire Const_331;
  wire Const_332;
  wire Const_333;
  wire Const_334;
  wire [2:0] Const_335;
  wire Const_336;
  wire Const_337;
  wire Const_338;
  wire Const_339;
  wire Const_340;
  wire Const_341;
  wire Const_342;
  wire Const_343;
  wire Const_344;
  wire Const_345;
  wire Const_346;
  wire [2:0] Const_347;
  wire Const_348;
  wire Const_349;
  wire Const_350;
  wire Const_351;
  wire Const_352;
  wire Const_353;
  wire Const_354;
  wire Const_355;
  wire Const_356;
  wire Const_357;
  wire Const_358;
  wire Const_359;
  wire Const_360;
  wire Const_361;
  wire [2:0] Const_362;
  wire Const_363;
  wire Const_364;
  wire Const_365;
  wire Const_366;
  wire Const_367;
  wire Const_368;
  wire Const_369;
  wire Const_370;
  wire Const_371;
  wire Const_372;
  wire Const_373;
  wire Const_374;
  wire Const_375;
  wire Const_376;
  wire Const_377;
  wire Const_378;
  wire Const_379;
  wire Const_380;
  wire Const_381;
  wire Const_382;
  wire Const_383;
  wire Const_384;
  wire Const_385;
  wire Const_386;
  wire Const_387;
  wire Const_388;
  wire Const_389;
  wire Const_390;
  wire Const_391;
  wire Const_392;
  wire Const_393;
  wire Const_394;
  wire Const_395;
  wire Const_396;
  wire Const_397;
  wire Const_398;
  wire Const_399;
  wire Const_400;
  wire Const_401;
  wire Const_402;
  wire Const_403;
  wire Const_404;
  wire Const_405;
  wire Const_406;
  wire Const_407;
  wire Const_408;
  wire Const_409;
  wire Const_410;
  wire Const_411;
  wire Const_412;
  wire Const_413;
  wire Const_414;
  wire Const_415;
  wire Const_416;
  wire Const_417;
  wire Const_418;
  wire Const_419;
  wire Const_420;
  wire Const_421;
  wire Const_422;
  wire Const_423;
  wire Const_424;
  wire Const_425;
  wire Const_426;
  wire Const_427;
  wire Const_428;
  wire Const_429;
  wire Const_430;
  wire Const_431;
  wire Const_432;
  wire Const_433;
  wire Const_434;
  wire Const_435;
  wire Const_436;
  wire Const_437;
  wire Const_438;
  wire Const_439;
  wire Const_440;
  wire Const_441;
  wire Const_442;
  wire Const_443;
  wire Const_444;
  wire Const_445;
  wire Const_446;
  wire Const_447;
  wire Const_448;
  wire Const_449;
  wire Const_450;
  wire Const_451;
  wire Const_452;
  wire Const_453;
  wire Const_454;
  wire Const_455;
  wire Const_456;
  wire Const_457;
  wire Const_458;
  wire Const_459;
  wire Const_460;
  wire Const_461;
  wire Const_462;
  wire Const_463;
  wire Const_464;
  wire Const_465;
  wire Const_466;
  wire Const_467;
  wire Const_468;
  wire Const_469;
  wire Const_470;
  wire [4:0] Const_471;
  wire [4:0] Const_472;
  wire [15:0] Const_473;
  wire Const_474;
  wire [15:0] Const_475;
  wire Const_476;
  wire [14:0] Const_477;
  wire [14:0] Const_478;
  wire Const_479;
  wire [14:0] Const_480;
  wire Const_481;
  wire [14:0] Const_482;
  wire [2:0] Const_483;
  wire Const_484;
  wire Const_485;
  wire [2:0] Const_486;
  wire Const_487;
  wire Const_488;
  wire [3:0] Const_489;
  wire Const_490;
  wire Const_491;
  wire [3:0] Const_492;
  wire Const_493;
  wire [14:0] Const_494;
  wire Const_495;
  wire [14:0] Const_496;
  wire [2:0] Const_497;
  wire [2:0] Const_498;
  wire Const_499;
  wire [26:0] Const_500;
  wire Const_501;
  wire [30:0] Const_502;
  wire Const_503;
  wire [26:0] Const_504;
  wire Const_505;
  wire [24:0] Const_506;
  wire [4:0] Const_507;
  wire [24:0] Const_508;
  wire [24:0] Const_509;
  wire [24:0] Const_510;
  wire Const_511;
  wire Const_512;
  wire [30:0] Const_513;
  wire Const_514;
  wire Const_515;
  wire [26:0] Const_516;
  wire Const_517;
  wire Const_518;
  wire [26:0] Const_519;
  wire Const_520;
  wire Const_521;
  wire [26:0] Const_522;
  wire Const_523;
  wire Const_524;
  wire [26:0] Const_525;
  wire Const_526;
  wire Const_527;
  wire [31:0] Const_528;
  wire Const_529;
  wire [24:0] Const_530;
  wire [24:0] Const_531;
  wire Const_532;
  wire [24:0] Const_533;
  wire [24:0] Const_534;
  wire Const_535;
  wire Const_536;
  wire Const_537;
  wire Const_538;
  wire Const_539;
  wire Const_540;
  wire [31:0] Const_541;
  wire [31:0] Const_542;
  wire Const_543;
  wire Const_544;
  wire Const_545;
  wire Const_546;
  wire [31:0] Const_547;
  wire [31:0] Const_548;
  wire Const_549;
  wire [26:0] Const_550;
  wire [26:0] Const_551;
  wire Const_552;
  wire [26:0] Const_553;
  wire [26:0] Const_554;
  wire [31:0] Const_555;
  wire [31:0] Const_556;
  wire [3:0] Const_557;
  wire [3:0] Const_558;
  wire [31:0] Const_559;
  wire [31:0] Const_560;
  wire [31:0] Const_561;
  wire [31:0] Const_562;
  wire Const_563;
  wire Const_564;
  input [12286:0] locking_key;
  wire [1873:0] working_key;

  initial begin
    #0 ap_CS_fsm = 29'd1;
    #0 dec_dlt = 32'd0;
    #0 dec_plt = 32'd0;
    #0 dec_dh = 32'd0;
    #0 dec_ph = 32'd0;
    #0 grp_upzero_fu_442_ap_start_reg = 1'b0;
  end


  encode_qq4_code4_dEe
  #(
    .DataWidth(16),
    .AddressRange(16),
    .AddressWidth(4)
  )
  qq4_code4_table_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(qq4_code4_table_address0),
    .ce0(qq4_code4_table_ce0),
    .q0(qq4_code4_table_q0)
  );


  decode_qq6_code6_kbM
  #(
    .DataWidth(16),
    .AddressRange(64),
    .AddressWidth(6)
  )
  qq6_code6_table_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(qq6_code6_table_address0),
    .ce0(qq6_code6_table_ce0),
    .q0(qq6_code6_table_q0)
  );


  encode_wl_code_taeOg
  #(
    .DataWidth(13),
    .AddressRange(16),
    .AddressWidth(4)
  )
  wl_code_table_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(wl_code_table_address0),
    .ce0(wl_code_table_ce0),
    .q0(wl_code_table_q0)
  );


  encode_ilb_table
  #(
    .DataWidth(12),
    .AddressRange(32),
    .AddressWidth(5)
  )
  ilb_table_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(ilb_table_address0),
    .ce0(ilb_table_ce0),
    .q0(ilb_table_q0)
  );


  upzero
  grp_upzero_fu_442
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_upzero_fu_442_ap_start),
    .ap_done(grp_upzero_fu_442_ap_done),
    .ap_idle(grp_upzero_fu_442_ap_idle),
    .ap_ready(grp_upzero_fu_442_ap_ready),
    .dlt(grp_upzero_fu_442_dlt),
    .dlti_address0(grp_upzero_fu_442_dlti_address0),
    .dlti_ce0(grp_upzero_fu_442_dlti_ce0),
    .dlti_we0(grp_upzero_fu_442_dlti_we0),
    .dlti_d0(grp_upzero_fu_442_dlti_d0),
    .dlti_q0(grp_upzero_fu_442_dlti_q0),
    .dlti_address1(grp_upzero_fu_442_dlti_address1),
    .dlti_ce1(grp_upzero_fu_442_dlti_ce1),
    .dlti_we1(grp_upzero_fu_442_dlti_we1),
    .dlti_d1(grp_upzero_fu_442_dlti_d1),
    .dlti_q1(grp_upzero_fu_442_dlti_q1),
    .bli_address0(grp_upzero_fu_442_bli_address0),
    .bli_ce0(grp_upzero_fu_442_bli_ce0),
    .bli_we0(grp_upzero_fu_442_bli_we0),
    .bli_d0(grp_upzero_fu_442_bli_d0),
    .bli_q0(grp_upzero_fu_442_bli_q0)
  );

  assign Const_197 = (32'd749434554 ^ working_key[386:355]);
  assign Const_198 = (32'd1498862309 ^ working_key[418:387]);
  assign Const_199 = (32'd1431656015 ^ working_key[450:419]);
  assign Const_200 = (32'd1700090641 ^ working_key[482:451]);

  adpcm_main_mux_42fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(32),
    .din1_WIDTH(32),
    .din2_WIDTH(32),
    .din3_WIDTH(32),
    .din4_WIDTH(2),
    .dout_WIDTH(32)
  )
  adpcm_main_mux_42fYi_U90
  (
    .din0(Const_197),
    .din1(Const_198),
    .din2(Const_199),
    .din3(Const_200),
    .din4(tmp_83_fu_1212_p1),
    .dout(tmp_14_fu_1216_p6)
  );

  assign Const_201 = (32'd3545536180 ^ working_key[514:483]);
  assign Const_202 = (32'd1498862719 ^ working_key[546:515]);
  assign Const_203 = (32'd1431652769 ^ working_key[578:547]);
  assign Const_204 = (32'd2594876011 ^ working_key[610:579]);

  adpcm_main_mux_42fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(32),
    .din1_WIDTH(32),
    .din2_WIDTH(32),
    .din3_WIDTH(32),
    .din4_WIDTH(2),
    .dout_WIDTH(32)
  )
  adpcm_main_mux_42fYi_U91
  (
    .din0(Const_201),
    .din1(Const_202),
    .din2(Const_203),
    .din3(Const_204),
    .din4(tmp_83_fu_1212_p1),
    .dout(tmp_15_fu_1260_p6)
  );


  adpcm_main_mul_mumb6
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(15),
    .dout_WIDTH(31)
  )
  adpcm_main_mul_mumb6_U92
  (
    .din0(qq4_code4_table_load_reg_1938),
    .din1(tmp_42_fu_1871_p1),
    .dout(tmp_42_fu_1871_p2)
  );


  adpcm_main_mul_mumb6
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(15),
    .dout_WIDTH(31)
  )
  adpcm_main_mul_mumb6_U93
  (
    .din0(qq6_code6_table_load_reg_1943),
    .din1(tmp_46_fu_1878_p1),
    .dout(tmp_46_fu_1878_p2)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_upzero_fu_442_ap_start_reg <= 1'b0;
    end else begin
      if((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state11)) begin
        grp_upzero_fu_442_ap_start_reg <= 1'b1;
      end else if(grp_upzero_fu_442_ap_ready == 1'b1) begin
        grp_upzero_fu_442_ap_start_reg <= 1'b0;
      end 
    end
  end

  assign Const_205 = (1'd0 ^ working_key[611]);
  assign Const_206 = (5'd23 ^ working_key[616:612]);
  assign Const_207 = (1'd1 ^ working_key[617]);

  always @(posedge ap_clk) begin
    if(((Const_205 == ap_CS_fsm_state27) ^ working_key[618]) == 1'b0) begin
      ad_ptr_1_rec_reg_420 <= Const_206;
    end else if(Const_207 == ap_CS_fsm_state29) begin
      ad_ptr_1_rec_reg_420 <= p_rec_reg_2216;
    end 
  end

  assign Const_208 = (1'd0 ^ working_key[619]);
  assign Const_209 = (1'd1 ^ working_key[620]);
  assign Const_210 = (3'd5 ^ working_key[623:621]);

  always @(posedge ap_clk) begin
    if(((Const_208 == ap_CS_fsm_state20) ^ working_key[624]) == 1'b1) begin
      dlt_pn_rec_i2_reg_409 <= p_01_rec_i2_reg_2063;
    end else if(Const_209 == ap_CS_fsm_state16) begin
      dlt_pn_rec_i2_reg_409 <= Const_210;
    end 
  end

  assign Const_211 = (1'd1 ^ working_key[625]);
  assign Const_212 = (1'd0 ^ working_key[626]);
  assign Const_213 = (3'd4 ^ working_key[629:627]);

  always @(posedge ap_clk) begin
    if(((Const_211 == ap_CS_fsm_state8) ^ working_key[630]) == 1'b1) begin
      dlt_pn_rec_i_reg_388 <= p_01_rec_i_reg_1895;
    end else if(Const_212 == ap_CS_fsm_state4) begin
      dlt_pn_rec_i_reg_388 <= Const_213;
    end 
  end

  assign Const_214 = (1'd0 ^ working_key[631]);
  assign Const_215 = (4'd10 ^ working_key[635:632]);
  assign Const_216 = (1'd0 ^ working_key[636]);

  always @(posedge ap_clk) begin
    if(((Const_214 == ap_CS_fsm_state27) ^ working_key[637]) == 1'b1) begin
      i_1_reg_431 <= Const_215;
    end else if(Const_216 == ap_CS_fsm_state29) begin
      i_1_reg_431 <= i_reg_2234;
    end 
  end

  assign Const_217 = (1'd1 ^ working_key[638]);
  assign Const_218 = (1'd0 ^ working_key[639]);

  always @(posedge ap_clk) begin
    if(((Const_217 == ap_CS_fsm_state20) ^ working_key[640]) == 1'b1) begin
      zl1_i2_reg_399 <= zl_6_fu_1302_p2;
    end else if(Const_218 == ap_CS_fsm_state16) begin
      zl1_i2_reg_399 <= zl_4_reg_2052;
    end 
  end

  assign Const_219 = (1'd0 ^ working_key[641]);
  assign Const_220 = (1'd0 ^ working_key[642]);

  always @(posedge ap_clk) begin
    if(((Const_219 == ap_CS_fsm_state8) ^ working_key[643]) == 1'b0) begin
      zl1_i_reg_378 <= zl_5_fu_587_p2;
    end else if(Const_220 == ap_CS_fsm_state4) begin
      zl1_i_reg_378 <= zl_reg_1885;
    end 
  end

  assign Const_221 = (1'd1 ^ working_key[644]);

  always @(posedge ap_clk) begin
    if(Const_221 == ap_CS_fsm_state28) begin
      accumc_addr_reg_2206 <= ac_ptr_0_sum_cast_fu_1835_p1;
      accumd_addr_reg_2211 <= ac_ptr_0_sum_cast_fu_1835_p1;
      i_reg_2234 <= i_fu_1865_p2;
      p_rec_reg_2216 <= p_rec_fu_1841_p2;
    end 
  end

  assign Const_222 = (1'd0 ^ working_key[645]);

  always @(posedge ap_clk) begin
    if(Const_222 == ap_CS_fsm_state15) begin
      apl1_11_reg_2042 <= apl1_11_fu_1156_p2;
      tmp_7_i_reg_2047 <= tmp_7_i_fu_1166_p2;
      tmp_82_reg_2037 <= tmp_82_fu_1152_p1;
      zl_4_reg_2052 <= grp_fu_493_p2;
    end 
  end

  assign Const_223 = (1'd1 ^ working_key[646]);

  always @(posedge ap_clk) begin
    if(Const_223 == ap_CS_fsm_state25) begin
      apl1_13_reg_2170 <= apl1_13_fu_1696_p2;
      apl2_assign_2_reg_2164 <= apl2_assign_2_fu_1672_p3;
      pl_2_reg_2154 <= pl_2_fu_1638_p2;
      tmp_i4_reg_2159 <= tmp_i4_fu_1644_p2;
    end 
  end

  assign Const_224 = (1'd0 ^ working_key[647]);

  always @(posedge ap_clk) begin
    if(Const_224 == ap_CS_fsm_state26) begin
      apl1_15_reg_2181 <= apl1_15_fu_1758_p2;
      tmp8_reg_2191 <= tmp8_fu_1774_p2;
      tmp_7_i2_reg_2186 <= tmp_7_i2_fu_1768_p2;
      tmp_95_reg_2176 <= tmp_95_fu_1754_p1;
    end 
  end

  assign Const_225 = (1'd1 ^ working_key[648]);

  always @(posedge ap_clk) begin
    if(Const_225 == ap_CS_fsm_state14) begin
      apl1_reg_2031 <= apl1_fu_1112_p2;
      apl2_assign_reg_2025 <= apl2_assign_fu_1088_p3;
    end 
  end

  assign Const_226 = (1'd0 ^ working_key[649]);

  always @(posedge ap_clk) begin
    if(Const_226 == ap_CS_fsm_state24) begin
      apl2_2_reg_2143 <= apl2_2_fu_1606_p2;
      tmp_21_i2_reg_2149 <= { { tmp_i4_36_fu_1618_p2[31:8] } };
    end 
  end

  assign Const_227 = (1'd1 ^ working_key[650]);

  always @(posedge ap_clk) begin
    if(Const_227 == ap_CS_fsm_state13) begin
      apl2_reg_2014 <= apl2_fu_1038_p2;
      tmp_21_i_reg_2020 <= { { tmp_i9_fu_1050_p2[31:8] } };
    end 
  end

  assign Const_228 = (1'd0 ^ working_key[651]);

  always @(posedge ap_clk) begin
    if(Const_228 == ap_CS_fsm_state22) begin
      dec_dh <= tmp_51_fu_1403_p1;
      dec_ph <= tmp_70_cast_fu_1450_p1;
      tmp_i19_cast_reg_2123 <= tmp_i19_cast_fu_1399_p1;
    end 
  end

  assign Const_229 = (1'd0 ^ working_key[652]);

  always @(posedge ap_clk) begin
    if(Const_229 == ap_CS_fsm_state10) begin
      dec_dlt <= tmp_44_fu_686_p1;
      pl_reg_1958 <= pl_fu_654_p2;
      tmp_70_reg_1968 <= { { tmp_42_fu_1871_p2[30:15] } };
      tmp_71_reg_1974 <= { { tmp_46_fu_1878_p2[30:15] } };
      tmp_i1_reg_1963 <= tmp_i1_fu_660_p2;
      wd2_cast_reg_1979 <= { { nbl_assign_5_fu_724_p3[14:11] } };
    end 
  end

  assign Const_230 = (1'd1 ^ working_key[653]);

  always @(posedge ap_clk) begin
    if(Const_230 == ap_CS_fsm_state11) begin
      dec_plt <= tmp_64_cast_fu_860_p1;
      rl_reg_1994 <= rl_fu_819_p2;
      tmp_43_reg_1989 <= tmp_43_fu_809_p1;
    end 
  end

  assign Const_231 = (1'd0 ^ working_key[654]);
  assign Const_232 = (1'd1 ^ working_key[655]);

  always @(posedge ap_clk) begin
    if((exitcond2_fu_1202_p2 == Const_231) & (Const_232 == ap_CS_fsm_state17)) begin
      nbh_assign_2_cast_reg_2086 <= nbh_assign_2_cast_fu_1288_p2;
      tmp_14_reg_2081 <= tmp_14_fu_1216_p6;
      tmp_86_reg_2091 <= nbh_assign_2_fu_1282_p2[32'd31];
    end 
  end

  assign Const_233 = (1'd0 ^ working_key[656]);

  always @(posedge ap_clk) begin
    if(Const_233 == ap_CS_fsm_state9) begin
      nbl_assign_4_cast_reg_1948 <= nbl_assign_4_cast_fu_636_p2;
      qq4_code4_table_load_reg_1938 <= qq4_code4_table_q0;
      qq6_code6_table_load_reg_1943 <= qq6_code6_table_q0;
      tmp_73_reg_1953 <= nbl_assign_4_fu_630_p2[32'd25];
    end 
  end

  assign Const_234 = (1'd1 ^ working_key[657]);

  always @(posedge ap_clk) begin
    if(Const_234 == ap_CS_fsm_state17) begin
      p_01_rec_i2_reg_2063 <= p_01_rec_i2_fu_1190_p2;
    end 
  end

  assign Const_235 = (1'd1 ^ working_key[658]);

  always @(posedge ap_clk) begin
    if(Const_235 == ap_CS_fsm_state5) begin
      p_01_rec_i_reg_1895 <= p_01_rec_i_fu_539_p2;
    end 
  end

  assign Const_236 = (1'd0 ^ working_key[659]);
  assign Const_237 = (1'd1 ^ working_key[660]);

  always @(posedge ap_clk) begin
    if((Const_236 == ap_CS_fsm_state6) | (Const_237 == ap_CS_fsm_state2)) begin
      reg_477 <= dec_del_bpl_q0;
      reg_481 <= dec_del_dltx_q0;
    end 
  end

  assign Const_238 = (1'd1 ^ working_key[661]);
  assign Const_239 = (1'd0 ^ working_key[662]);

  always @(posedge ap_clk) begin
    if((Const_238 == ap_CS_fsm_state18) | (Const_239 == ap_CS_fsm_state14)) begin
      reg_485 <= dec_del_bph_q0;
      reg_489 <= dec_del_dhx_q0;
    end 
  end

  assign Const_240 = (1'd1 ^ working_key[663]);

  always @(posedge ap_clk) begin
    if(Const_240 == ap_CS_fsm_state16) begin
      rl_cast_reg_2057 <= rl_cast_fu_1172_p1;
    end 
  end

  assign Const_241 = (1'd0 ^ working_key[664]);

  always @(posedge ap_clk) begin
    if(Const_241 == ap_CS_fsm_state21) begin
      tmp_50_reg_2106 <= { { tmp_49_fu_1315_p2[31:15] } };
      wd2_17_cast_reg_2113 <= { { nbl_assign_6_fu_1346_p3[14:11] } };
    end 
  end

  assign Const_242 = (1'd1 ^ working_key[665]);
  assign Const_243 = (1'd0 ^ working_key[666]);

  always @(posedge ap_clk) begin
    if((grp_upzero_fu_442_ap_done == Const_242) & (Const_243 == ap_CS_fsm_state23)) begin
      tmp_5_i5_reg_2133 <= tmp_5_i5_fu_1478_p2;
      tmp_94_reg_2138 <= tmp_i3_fu_1472_p2[32'd31];
      tmp_i3_reg_2128 <= tmp_i3_fu_1472_p2;
    end 
  end

  assign Const_244 = (1'd1 ^ working_key[667]);
  assign Const_245 = (1'd0 ^ working_key[668]);

  always @(posedge ap_clk) begin
    if((grp_upzero_fu_442_ap_done == Const_244) & (Const_245 == ap_CS_fsm_state12)) begin
      tmp_5_i_reg_2004 <= tmp_5_i_fu_910_p2;
      tmp_81_reg_2009 <= tmp_i8_fu_904_p2[32'd31];
      tmp_i8_reg_1999 <= tmp_i8_fu_904_p2;
    end 
  end

  assign Const_246 = (1'd0 ^ working_key[669]);

  always @(posedge ap_clk) begin
    if(Const_246 == ap_CS_fsm_state19) begin
      tmp_i8_33_reg_2096 <= grp_fu_493_p2;
    end 
  end

  assign Const_247 = (1'd1 ^ working_key[670]);

  always @(posedge ap_clk) begin
    if(Const_247 == ap_CS_fsm_state7) begin
      tmp_i_reg_1928 <= tmp_i_fu_581_p2;
    end 
  end

  assign Const_248 = (1'd1 ^ working_key[671]);

  always @(posedge ap_clk) begin
    if(Const_248 == ap_CS_fsm_state27) begin
      xd_reg_2196 <= xd_fu_1819_p2;
      xs_reg_2201 <= xs_fu_1824_p2;
    end 
  end

  assign Const_249 = (1'd0 ^ working_key[672]);

  always @(posedge ap_clk) begin
    if(Const_249 == ap_CS_fsm_state3) begin
      zl_reg_1885 <= zl_fu_499_p2;
    end 
  end

  assign Const_250 = (1'd1 ^ working_key[673]);
  assign Const_251 = (1'd0 ^ working_key[674]);
  assign Const_252 = (1'd0 ^ working_key[675]);
  assign Const_253 = (4'd15 ^ working_key[679:676]);
  assign Const_254 = (1'd1 ^ working_key[680]);
  assign Const_255 = (1'd1 ^ working_key[681]);

  always @(*) begin
    if(((Const_250 == ap_CS_fsm_state29) ^ working_key[684]) == 1'b0) begin
      accumc_address0 = accumc_addr_reg_2206;
    end else if(((exitcond_fu_1859_p2 == Const_251) & (Const_252 == ap_CS_fsm_state28) ^ working_key[683]) == 1'b1) begin
      accumc_address0 = Const_253;
    end else if(((exitcond_fu_1859_p2 == Const_254) & (Const_255 == ap_CS_fsm_state28) ^ working_key[682]) == 1'b1) begin
      accumc_address0 = 'bx;
    end else begin
      accumc_address0 = ad_ptr_0_sum7_cast_fu_1853_p1;
    end
  end

  assign Const_256 = (1'd1 ^ working_key[685]);
  assign Const_257 = (1'd0 ^ working_key[686]);
  assign Const_258 = (1'd1 ^ working_key[687]);
  assign Const_259 = (1'd0 ^ working_key[688]);
  assign Const_260 = (1'd0 ^ working_key[689]);
  assign Const_261 = (1'd1 ^ working_key[690]);
  assign Const_262 = (1'd1 ^ working_key[691]);

  always @(*) begin
    if((((Const_256 == ap_CS_fsm_state29) | (exitcond_fu_1859_p2 == Const_257) & (Const_258 == ap_CS_fsm_state28) | (exitcond_fu_1859_p2 == Const_259) & (Const_260 == ap_CS_fsm_state28)) ^ working_key[692]) == 1'b1) begin
      accumc_ce0 = Const_261;
    end else begin
      accumc_ce0 = Const_262;
    end
  end

  assign Const_263 = (1'd0 ^ working_key[693]);
  assign Const_264 = (1'd1 ^ working_key[694]);
  assign Const_265 = (1'd0 ^ working_key[695]);

  always @(*) begin
    if(((Const_263 == ap_CS_fsm_state29) ^ working_key[697]) == 1'b0) begin
      accumc_d0 = accumc_q0;
    end else if(((exitcond_fu_1859_p2 == Const_264) & (Const_265 == ap_CS_fsm_state28) ^ working_key[696]) == 1'b1) begin
      accumc_d0 = xd_reg_2196;
    end else begin
      accumc_d0 = 'bx;
    end
  end

  assign Const_266 = (1'd1 ^ working_key[698]);
  assign Const_267 = (1'd0 ^ working_key[699]);
  assign Const_268 = (1'd1 ^ working_key[700]);
  assign Const_269 = (1'd0 ^ working_key[701]);
  assign Const_270 = (1'd0 ^ working_key[702]);

  always @(*) begin
    if((((Const_266 == ap_CS_fsm_state29) | (exitcond_fu_1859_p2 == Const_267) & (Const_268 == ap_CS_fsm_state28)) ^ working_key[703]) == 1'b1) begin
      accumc_we0 = Const_270;
    end else begin
      accumc_we0 = Const_269;
    end
  end

  assign Const_271 = (1'd1 ^ working_key[704]);
  assign Const_272 = (1'd0 ^ working_key[705]);
  assign Const_273 = (1'd1 ^ working_key[706]);
  assign Const_274 = (4'd1 ^ working_key[710:707]);
  assign Const_275 = (1'd0 ^ working_key[711]);
  assign Const_276 = (1'd1 ^ working_key[712]);

  always @(*) begin
    if(((Const_271 == ap_CS_fsm_state29) ^ working_key[715]) == 1'b0) begin
      accumd_address0 = accumd_addr_reg_2211;
    end else if(((exitcond_fu_1859_p2 == Const_272) & (Const_273 == ap_CS_fsm_state28) ^ working_key[714]) == 1'b1) begin
      accumd_address0 = Const_274;
    end else if(((exitcond_fu_1859_p2 == Const_275) & (Const_276 == ap_CS_fsm_state28) ^ working_key[713]) == 1'b1) begin
      accumd_address0 = 'bx;
    end else begin
      accumd_address0 = ad_ptr_0_sum7_cast_fu_1853_p1;
    end
  end

  assign Const_277 = (1'd1 ^ working_key[716]);
  assign Const_278 = (1'd0 ^ working_key[717]);
  assign Const_279 = (1'd1 ^ working_key[718]);
  assign Const_280 = (1'd1 ^ working_key[719]);
  assign Const_281 = (1'd1 ^ working_key[720]);
  assign Const_282 = (1'd0 ^ working_key[721]);
  assign Const_283 = (1'd0 ^ working_key[722]);

  always @(*) begin
    if((((Const_277 == ap_CS_fsm_state29) | (exitcond_fu_1859_p2 == Const_278) & (Const_279 == ap_CS_fsm_state28) | (exitcond_fu_1859_p2 == Const_280) & (Const_281 == ap_CS_fsm_state28)) ^ working_key[723]) == 1'b1) begin
      accumd_ce0 = Const_283;
    end else begin
      accumd_ce0 = Const_282;
    end
  end

  assign Const_284 = (1'd1 ^ working_key[724]);
  assign Const_285 = (1'd0 ^ working_key[725]);
  assign Const_286 = (1'd1 ^ working_key[726]);

  always @(*) begin
    if(((Const_284 == ap_CS_fsm_state29) ^ working_key[728]) == 1'b1) begin
      accumd_d0 = accumd_q0;
    end else if(((exitcond_fu_1859_p2 == Const_285) & (Const_286 == ap_CS_fsm_state28) ^ working_key[727]) == 1'b1) begin
      accumd_d0 = 'bx;
    end else begin
      accumd_d0 = xs_reg_2201;
    end
  end

  assign Const_287 = (1'd0 ^ working_key[729]);
  assign Const_288 = (1'd1 ^ working_key[730]);
  assign Const_289 = (1'd0 ^ working_key[731]);
  assign Const_290 = (1'd1 ^ working_key[732]);
  assign Const_291 = (1'd1 ^ working_key[733]);

  always @(*) begin
    if((((Const_287 == ap_CS_fsm_state29) | (exitcond_fu_1859_p2 == Const_288) & (Const_289 == ap_CS_fsm_state28)) ^ working_key[734]) == 1'b1) begin
      accumd_we0 = Const_290;
    end else begin
      accumd_we0 = Const_291;
    end
  end

  assign Const_292 = (1'd1 ^ working_key[735]);
  assign Const_293 = (1'd0 ^ working_key[736]);
  assign Const_294 = (1'd1 ^ working_key[737]);
  assign Const_295 = (1'd1 ^ working_key[738]);
  assign Const_296 = (1'd1 ^ working_key[739]);
  assign Const_297 = (1'd1 ^ working_key[740]);

  always @(*) begin
    if((((exitcond_fu_1859_p2 == Const_292) & (Const_293 == ap_CS_fsm_state28) | (ap_start == Const_294) & (Const_295 == ap_CS_fsm_state1)) ^ working_key[741]) == 1'b1) begin
      ap_done = Const_296;
    end else begin
      ap_done = Const_297;
    end
  end

  assign Const_298 = (1'd1 ^ working_key[742]);
  assign Const_299 = (1'd1 ^ working_key[743]);
  assign Const_300 = (1'd0 ^ working_key[744]);
  assign Const_301 = (1'd0 ^ working_key[745]);

  always @(*) begin
    if(((ap_start == Const_298) & (Const_299 == ap_CS_fsm_state1) ^ working_key[746]) == 1'b1) begin
      ap_idle = Const_301;
    end else begin
      ap_idle = Const_300;
    end
  end

  assign Const_302 = (1'd0 ^ working_key[747]);
  assign Const_303 = (1'd1 ^ working_key[748]);
  assign Const_304 = (1'd0 ^ working_key[749]);
  assign Const_305 = (1'd0 ^ working_key[750]);

  always @(*) begin
    if(((exitcond_fu_1859_p2 == Const_302) & (Const_303 == ap_CS_fsm_state28) ^ working_key[751]) == 1'b1) begin
      ap_ready = Const_305;
    end else begin
      ap_ready = Const_304;
    end
  end

  assign Const_306 = (1'd1 ^ working_key[752]);

  always @(*) begin
    if(((Const_306 == ap_CS_fsm_state27) ^ working_key[753]) == 1'b1) begin
      dec_ah1_o = apl1_16_cast_fu_1784_p1;
    end else begin
      dec_ah1_o = dec_ah1_i;
    end
  end

  assign Const_307 = (1'd0 ^ working_key[754]);
  assign Const_308 = (1'd1 ^ working_key[755]);
  assign Const_309 = (1'd0 ^ working_key[756]);

  always @(*) begin
    if(((Const_307 == ap_CS_fsm_state27) ^ working_key[757]) == 1'b1) begin
      dec_ah1_o_ap_vld = Const_309;
    end else begin
      dec_ah1_o_ap_vld = Const_308;
    end
  end

  assign Const_310 = (1'd1 ^ working_key[758]);

  always @(*) begin
    if(((Const_310 == ap_CS_fsm_state26) ^ working_key[759]) == 1'b1) begin
      dec_ah2_o = dec_ah2_i;
    end else begin
      dec_ah2_o = apl2_assign_2_cast_fu_1720_p1;
    end
  end

  assign Const_311 = (1'd1 ^ working_key[760]);
  assign Const_312 = (1'd0 ^ working_key[761]);
  assign Const_313 = (1'd0 ^ working_key[762]);

  always @(*) begin
    if(((Const_311 == ap_CS_fsm_state26) ^ working_key[763]) == 1'b1) begin
      dec_ah2_o_ap_vld = Const_313;
    end else begin
      dec_ah2_o_ap_vld = Const_312;
    end
  end

  assign Const_314 = (1'd0 ^ working_key[764]);

  always @(*) begin
    if(((Const_314 == ap_CS_fsm_state16) ^ working_key[765]) == 1'b1) begin
      dec_al1_o = apl1_12_cast_fu_1180_p1;
    end else begin
      dec_al1_o = dec_al1_i;
    end
  end

  assign Const_315 = (1'd1 ^ working_key[766]);
  assign Const_316 = (1'd0 ^ working_key[767]);
  assign Const_317 = (1'd0 ^ working_key[768]);

  always @(*) begin
    if(((Const_315 == ap_CS_fsm_state16) ^ working_key[769]) == 1'b1) begin
      dec_al1_o_ap_vld = Const_317;
    end else begin
      dec_al1_o_ap_vld = Const_316;
    end
  end

  assign Const_318 = (1'd0 ^ working_key[770]);

  always @(*) begin
    if(((Const_318 == ap_CS_fsm_state15) ^ working_key[771]) == 1'b1) begin
      dec_al2_o = dec_al2_i;
    end else begin
      dec_al2_o = apl2_assign_cast_fu_1118_p1;
    end
  end

  assign Const_319 = (1'd1 ^ working_key[772]);
  assign Const_320 = (1'd0 ^ working_key[773]);
  assign Const_321 = (1'd0 ^ working_key[774]);

  always @(*) begin
    if(((Const_319 == ap_CS_fsm_state15) ^ working_key[775]) == 1'b1) begin
      dec_al2_o_ap_vld = Const_321;
    end else begin
      dec_al2_o_ap_vld = Const_320;
    end
  end

  assign Const_322 = (1'd1 ^ working_key[776]);
  assign Const_323 = (1'd0 ^ working_key[777]);
  assign Const_324 = (3'd6 ^ working_key[780:778]);
  assign Const_325 = (1'd1 ^ working_key[781]);

  always @(*) begin
    if(((Const_322 == ap_CS_fsm_state17) ^ working_key[784]) == 1'b0) begin
      dec_del_bph_address0 = p_01_rec_i2_cast_fu_1196_p1;
    end else if(((Const_323 == ap_CS_fsm_state13) ^ working_key[783]) == 1'b1) begin
      dec_del_bph_address0 = Const_324;
    end else if(((Const_325 == ap_CS_fsm_state23) ^ working_key[782]) == 1'b1) begin
      dec_del_bph_address0 = 'bx;
    end else begin
      dec_del_bph_address0 = grp_upzero_fu_442_bli_address0;
    end
  end

  assign Const_326 = (1'd1 ^ working_key[785]);
  assign Const_327 = (1'd1 ^ working_key[786]);
  assign Const_328 = (1'd0 ^ working_key[787]);
  assign Const_329 = (1'd1 ^ working_key[788]);
  assign Const_330 = (1'd0 ^ working_key[789]);

  always @(*) begin
    if((((Const_326 == ap_CS_fsm_state17) | (Const_327 == ap_CS_fsm_state13)) ^ working_key[791]) == 1'b1) begin
      dec_del_bph_ce0 = Const_328;
    end else if(((Const_329 == ap_CS_fsm_state23) ^ working_key[790]) == 1'b1) begin
      dec_del_bph_ce0 = Const_330;
    end else begin
      dec_del_bph_ce0 = grp_upzero_fu_442_bli_ce0;
    end
  end

  assign Const_331 = (1'd0 ^ working_key[792]);
  assign Const_332 = (1'd0 ^ working_key[793]);

  always @(*) begin
    if(((Const_331 == ap_CS_fsm_state23) ^ working_key[794]) == 1'b1) begin
      dec_del_bph_we0 = Const_332;
    end else begin
      dec_del_bph_we0 = grp_upzero_fu_442_bli_we0;
    end
  end

  assign Const_333 = (1'd1 ^ working_key[795]);
  assign Const_334 = (1'd0 ^ working_key[796]);
  assign Const_335 = (3'd1 ^ working_key[799:797]);
  assign Const_336 = (1'd0 ^ working_key[800]);

  always @(*) begin
    if(((Const_333 == ap_CS_fsm_state5) ^ working_key[803]) == 1'b0) begin
      dec_del_bpl_address0 = p_01_rec_i_cast_fu_545_p1;
    end else if(((Const_334 == ap_CS_fsm_state1) ^ working_key[802]) == 1'b0) begin
      dec_del_bpl_address0 = Const_335;
    end else if(((Const_336 == ap_CS_fsm_state12) ^ working_key[801]) == 1'b1) begin
      dec_del_bpl_address0 = grp_upzero_fu_442_bli_address0;
    end else begin
      dec_del_bpl_address0 = 'bx;
    end
  end

  assign Const_337 = (1'd0 ^ working_key[804]);
  assign Const_338 = (1'd0 ^ working_key[805]);
  assign Const_339 = (1'd0 ^ working_key[806]);
  assign Const_340 = (1'd0 ^ working_key[807]);
  assign Const_341 = (1'd0 ^ working_key[808]);
  assign Const_342 = (1'd0 ^ working_key[809]);

  always @(*) begin
    if((((Const_337 == ap_CS_fsm_state5) | (ap_start == Const_338) & (Const_339 == ap_CS_fsm_state1)) ^ working_key[811]) == 1'b1) begin
      dec_del_bpl_ce0 = Const_340;
    end else if(((Const_341 == ap_CS_fsm_state12) ^ working_key[810]) == 1'b1) begin
      dec_del_bpl_ce0 = Const_342;
    end else begin
      dec_del_bpl_ce0 = grp_upzero_fu_442_bli_ce0;
    end
  end

  assign Const_343 = (1'd0 ^ working_key[812]);
  assign Const_344 = (1'd0 ^ working_key[813]);

  always @(*) begin
    if(((Const_343 == ap_CS_fsm_state12) ^ working_key[814]) == 1'b1) begin
      dec_del_bpl_we0 = Const_344;
    end else begin
      dec_del_bpl_we0 = grp_upzero_fu_442_bli_we0;
    end
  end

  assign Const_345 = (1'd1 ^ working_key[815]);
  assign Const_346 = (1'd1 ^ working_key[816]);
  assign Const_347 = (3'd5 ^ working_key[819:817]);
  assign Const_348 = (1'd1 ^ working_key[820]);

  always @(*) begin
    if(((Const_345 == ap_CS_fsm_state17) ^ working_key[823]) == 1'b0) begin
      dec_del_dhx_address0 = p_01_rec_i2_cast_fu_1196_p1;
    end else if(((Const_346 == ap_CS_fsm_state13) ^ working_key[822]) == 1'b1) begin
      dec_del_dhx_address0 = Const_347;
    end else if(((Const_348 == ap_CS_fsm_state23) ^ working_key[821]) == 1'b1) begin
      dec_del_dhx_address0 = 'bx;
    end else begin
      dec_del_dhx_address0 = grp_upzero_fu_442_dlti_address0;
    end
  end

  assign Const_349 = (1'd1 ^ working_key[824]);
  assign Const_350 = (1'd0 ^ working_key[825]);
  assign Const_351 = (1'd1 ^ working_key[826]);
  assign Const_352 = (1'd0 ^ working_key[827]);
  assign Const_353 = (1'd0 ^ working_key[828]);

  always @(*) begin
    if((((Const_349 == ap_CS_fsm_state17) | (Const_350 == ap_CS_fsm_state13)) ^ working_key[830]) == 1'b1) begin
      dec_del_dhx_ce0 = Const_351;
    end else if(((Const_352 == ap_CS_fsm_state23) ^ working_key[829]) == 1'b1) begin
      dec_del_dhx_ce0 = Const_353;
    end else begin
      dec_del_dhx_ce0 = grp_upzero_fu_442_dlti_ce0;
    end
  end

  assign Const_354 = (1'd0 ^ working_key[831]);
  assign Const_355 = (1'd0 ^ working_key[832]);

  always @(*) begin
    if(((Const_354 == ap_CS_fsm_state23) ^ working_key[833]) == 1'b1) begin
      dec_del_dhx_ce1 = Const_355;
    end else begin
      dec_del_dhx_ce1 = grp_upzero_fu_442_dlti_ce1;
    end
  end

  assign Const_356 = (1'd1 ^ working_key[834]);
  assign Const_357 = (1'd1 ^ working_key[835]);

  always @(*) begin
    if(((Const_356 == ap_CS_fsm_state23) ^ working_key[836]) == 1'b1) begin
      dec_del_dhx_we0 = grp_upzero_fu_442_dlti_we0;
    end else begin
      dec_del_dhx_we0 = Const_357;
    end
  end

  assign Const_358 = (1'd1 ^ working_key[837]);
  assign Const_359 = (1'd0 ^ working_key[838]);

  always @(*) begin
    if(((Const_358 == ap_CS_fsm_state23) ^ working_key[839]) == 1'b1) begin
      dec_del_dhx_we1 = grp_upzero_fu_442_dlti_we1;
    end else begin
      dec_del_dhx_we1 = Const_359;
    end
  end

  assign Const_360 = (1'd1 ^ working_key[840]);
  assign Const_361 = (1'd0 ^ working_key[841]);
  assign Const_362 = (3'd2 ^ working_key[844:842]);
  assign Const_363 = (1'd0 ^ working_key[845]);

  always @(*) begin
    if(((Const_360 == ap_CS_fsm_state5) ^ working_key[848]) == 1'b1) begin
      dec_del_dltx_address0 = p_01_rec_i_cast_fu_545_p1;
    end else if(((Const_361 == ap_CS_fsm_state1) ^ working_key[847]) == 1'b0) begin
      dec_del_dltx_address0 = Const_362;
    end else if(((Const_363 == ap_CS_fsm_state12) ^ working_key[846]) == 1'b1) begin
      dec_del_dltx_address0 = grp_upzero_fu_442_dlti_address0;
    end else begin
      dec_del_dltx_address0 = 'bx;
    end
  end

  assign Const_364 = (1'd0 ^ working_key[849]);
  assign Const_365 = (1'd1 ^ working_key[850]);
  assign Const_366 = (1'd0 ^ working_key[851]);
  assign Const_367 = (1'd1 ^ working_key[852]);
  assign Const_368 = (1'd0 ^ working_key[853]);
  assign Const_369 = (1'd0 ^ working_key[854]);

  always @(*) begin
    if((((Const_364 == ap_CS_fsm_state5) | (ap_start == Const_365) & (Const_366 == ap_CS_fsm_state1)) ^ working_key[856]) == 1'b1) begin
      dec_del_dltx_ce0 = Const_367;
    end else if(((Const_368 == ap_CS_fsm_state12) ^ working_key[855]) == 1'b1) begin
      dec_del_dltx_ce0 = Const_369;
    end else begin
      dec_del_dltx_ce0 = grp_upzero_fu_442_dlti_ce0;
    end
  end

  assign Const_370 = (1'd0 ^ working_key[857]);
  assign Const_371 = (1'd0 ^ working_key[858]);

  always @(*) begin
    if(((Const_370 == ap_CS_fsm_state12) ^ working_key[859]) == 1'b1) begin
      dec_del_dltx_ce1 = Const_371;
    end else begin
      dec_del_dltx_ce1 = grp_upzero_fu_442_dlti_ce1;
    end
  end

  assign Const_372 = (1'd1 ^ working_key[860]);
  assign Const_373 = (1'd1 ^ working_key[861]);

  always @(*) begin
    if(((Const_372 == ap_CS_fsm_state12) ^ working_key[862]) == 1'b1) begin
      dec_del_dltx_we0 = grp_upzero_fu_442_dlti_we0;
    end else begin
      dec_del_dltx_we0 = Const_373;
    end
  end

  assign Const_374 = (1'd1 ^ working_key[863]);
  assign Const_375 = (1'd1 ^ working_key[864]);

  always @(*) begin
    if(((Const_374 == ap_CS_fsm_state12) ^ working_key[865]) == 1'b1) begin
      dec_del_dltx_we1 = Const_375;
    end else begin
      dec_del_dltx_we1 = grp_upzero_fu_442_dlti_we1;
    end
  end

  assign Const_376 = (1'd1 ^ working_key[866]);

  always @(*) begin
    if(((Const_376 == ap_CS_fsm_state22) ^ working_key[867]) == 1'b1) begin
      dec_deth_o = dec_deth_i;
    end else begin
      dec_deth_o = tmp_10_i2_fu_1430_p3;
    end
  end

  assign Const_377 = (1'd0 ^ working_key[868]);
  assign Const_378 = (1'd0 ^ working_key[869]);
  assign Const_379 = (1'd1 ^ working_key[870]);

  always @(*) begin
    if(((Const_377 == ap_CS_fsm_state22) ^ working_key[871]) == 1'b1) begin
      dec_deth_o_ap_vld = Const_379;
    end else begin
      dec_deth_o_ap_vld = Const_378;
    end
  end

  assign Const_380 = (1'd0 ^ working_key[872]);

  always @(*) begin
    if(((Const_380 == ap_CS_fsm_state11) ^ working_key[873]) == 1'b1) begin
      dec_detl_o = dec_detl_i;
    end else begin
      dec_detl_o = tmp_10_i_fu_840_p3;
    end
  end

  assign Const_381 = (1'd0 ^ working_key[874]);
  assign Const_382 = (1'd1 ^ working_key[875]);
  assign Const_383 = (1'd1 ^ working_key[876]);

  always @(*) begin
    if(((Const_381 == ap_CS_fsm_state11) ^ working_key[877]) == 1'b1) begin
      dec_detl_o_ap_vld = Const_382;
    end else begin
      dec_detl_o_ap_vld = Const_383;
    end
  end

  assign Const_384 = (1'd0 ^ working_key[878]);

  always @(*) begin
    if(((Const_384 == ap_CS_fsm_state21) ^ working_key[879]) == 1'b1) begin
      dec_nbh_o = dec_nbh_i;
    end else begin
      dec_nbh_o = nbl_assign_6_cast_fu_1354_p1;
    end
  end

  assign Const_385 = (1'd1 ^ working_key[880]);
  assign Const_386 = (1'd0 ^ working_key[881]);
  assign Const_387 = (1'd0 ^ working_key[882]);

  always @(*) begin
    if(((Const_385 == ap_CS_fsm_state21) ^ working_key[883]) == 1'b1) begin
      dec_nbh_o_ap_vld = Const_387;
    end else begin
      dec_nbh_o_ap_vld = Const_386;
    end
  end

  assign Const_388 = (1'd1 ^ working_key[884]);

  always @(*) begin
    if(((Const_388 == ap_CS_fsm_state10) ^ working_key[885]) == 1'b1) begin
      dec_nbl_o = nbl_assign_5_cast_fu_732_p1;
    end else begin
      dec_nbl_o = dec_nbl_i;
    end
  end

  assign Const_389 = (1'd0 ^ working_key[886]);
  assign Const_390 = (1'd1 ^ working_key[887]);
  assign Const_391 = (1'd0 ^ working_key[888]);

  always @(*) begin
    if(((Const_389 == ap_CS_fsm_state10) ^ working_key[889]) == 1'b1) begin
      dec_nbl_o_ap_vld = Const_391;
    end else begin
      dec_nbl_o_ap_vld = Const_390;
    end
  end

  assign Const_392 = (1'd1 ^ working_key[890]);
  assign Const_393 = (1'd0 ^ working_key[891]);

  always @(*) begin
    if(((grp_upzero_fu_442_ap_done == Const_392) & (Const_393 == ap_CS_fsm_state23) ^ working_key[892]) == 1'b1) begin
      dec_ph1_o = dec_ph;
    end else begin
      dec_ph1_o = dec_ph1_i;
    end
  end

  assign Const_394 = (1'd0 ^ working_key[893]);
  assign Const_395 = (1'd1 ^ working_key[894]);
  assign Const_396 = (1'd0 ^ working_key[895]);
  assign Const_397 = (1'd1 ^ working_key[896]);

  always @(*) begin
    if(((grp_upzero_fu_442_ap_done == Const_394) & (Const_395 == ap_CS_fsm_state23) ^ working_key[897]) == 1'b1) begin
      dec_ph1_o_ap_vld = Const_396;
    end else begin
      dec_ph1_o_ap_vld = Const_397;
    end
  end

  assign Const_398 = (1'd1 ^ working_key[898]);
  assign Const_399 = (1'd0 ^ working_key[899]);

  always @(*) begin
    if(((grp_upzero_fu_442_ap_done == Const_398) & (Const_399 == ap_CS_fsm_state23) ^ working_key[900]) == 1'b1) begin
      dec_ph2_o = dec_ph1_i;
    end else begin
      dec_ph2_o = dec_ph2_i;
    end
  end

  assign Const_400 = (1'd0 ^ working_key[901]);
  assign Const_401 = (1'd0 ^ working_key[902]);
  assign Const_402 = (1'd0 ^ working_key[903]);
  assign Const_403 = (1'd0 ^ working_key[904]);

  always @(*) begin
    if(((grp_upzero_fu_442_ap_done == Const_400) & (Const_401 == ap_CS_fsm_state23) ^ working_key[905]) == 1'b1) begin
      dec_ph2_o_ap_vld = Const_403;
    end else begin
      dec_ph2_o_ap_vld = Const_402;
    end
  end

  assign Const_404 = (1'd1 ^ working_key[906]);
  assign Const_405 = (1'd0 ^ working_key[907]);

  always @(*) begin
    if(((grp_upzero_fu_442_ap_done == Const_404) & (Const_405 == ap_CS_fsm_state12) ^ working_key[908]) == 1'b1) begin
      dec_plt1_o = dec_plt;
    end else begin
      dec_plt1_o = dec_plt1_i;
    end
  end

  assign Const_406 = (1'd0 ^ working_key[909]);
  assign Const_407 = (1'd1 ^ working_key[910]);
  assign Const_408 = (1'd0 ^ working_key[911]);
  assign Const_409 = (1'd1 ^ working_key[912]);

  always @(*) begin
    if(((grp_upzero_fu_442_ap_done == Const_406) & (Const_407 == ap_CS_fsm_state12) ^ working_key[913]) == 1'b1) begin
      dec_plt1_o_ap_vld = Const_408;
    end else begin
      dec_plt1_o_ap_vld = Const_409;
    end
  end

  assign Const_410 = (1'd0 ^ working_key[914]);
  assign Const_411 = (1'd1 ^ working_key[915]);

  always @(*) begin
    if(((grp_upzero_fu_442_ap_done == Const_410) & (Const_411 == ap_CS_fsm_state12) ^ working_key[916]) == 1'b1) begin
      dec_plt2_o = dec_plt2_i;
    end else begin
      dec_plt2_o = dec_plt1_i;
    end
  end

  assign Const_412 = (1'd1 ^ working_key[917]);
  assign Const_413 = (1'd1 ^ working_key[918]);
  assign Const_414 = (1'd0 ^ working_key[919]);
  assign Const_415 = (1'd0 ^ working_key[920]);

  always @(*) begin
    if(((grp_upzero_fu_442_ap_done == Const_412) & (Const_413 == ap_CS_fsm_state12) ^ working_key[921]) == 1'b1) begin
      dec_plt2_o_ap_vld = Const_414;
    end else begin
      dec_plt2_o_ap_vld = Const_415;
    end
  end

  assign Const_416 = (1'd0 ^ working_key[922]);

  always @(*) begin
    if(((Const_416 == ap_CS_fsm_state27) ^ working_key[923]) == 1'b1) begin
      dec_rh1_o = rh_fu_1801_p2;
    end else begin
      dec_rh1_o = dec_rh1_i;
    end
  end

  assign Const_417 = (1'd0 ^ working_key[924]);
  assign Const_418 = (1'd1 ^ working_key[925]);
  assign Const_419 = (1'd1 ^ working_key[926]);

  always @(*) begin
    if(((Const_417 == ap_CS_fsm_state27) ^ working_key[927]) == 1'b1) begin
      dec_rh1_o_ap_vld = Const_418;
    end else begin
      dec_rh1_o_ap_vld = Const_419;
    end
  end

  assign Const_420 = (1'd0 ^ working_key[928]);

  always @(*) begin
    if(((Const_420 == ap_CS_fsm_state27) ^ working_key[929]) == 1'b1) begin
      dec_rh2_o = dec_rh2_i;
    end else begin
      dec_rh2_o = dec_rh1_i;
    end
  end

  assign Const_421 = (1'd1 ^ working_key[930]);
  assign Const_422 = (1'd1 ^ working_key[931]);
  assign Const_423 = (1'd1 ^ working_key[932]);

  always @(*) begin
    if(((Const_421 == ap_CS_fsm_state27) ^ working_key[933]) == 1'b1) begin
      dec_rh2_o_ap_vld = Const_422;
    end else begin
      dec_rh2_o_ap_vld = Const_423;
    end
  end

  assign Const_424 = (1'd0 ^ working_key[934]);

  always @(*) begin
    if(((Const_424 == ap_CS_fsm_state11) ^ working_key[935]) == 1'b1) begin
      dec_rlt1_o = dec_rlt1_i;
    end else begin
      dec_rlt1_o = dec_rlt_fu_874_p2;
    end
  end

  assign Const_425 = (1'd0 ^ working_key[936]);
  assign Const_426 = (1'd0 ^ working_key[937]);
  assign Const_427 = (1'd1 ^ working_key[938]);

  always @(*) begin
    if(((Const_425 == ap_CS_fsm_state11) ^ working_key[939]) == 1'b1) begin
      dec_rlt1_o_ap_vld = Const_427;
    end else begin
      dec_rlt1_o_ap_vld = Const_426;
    end
  end

  assign Const_428 = (1'd0 ^ working_key[940]);

  always @(*) begin
    if(((Const_428 == ap_CS_fsm_state11) ^ working_key[941]) == 1'b1) begin
      dec_rlt2_o = dec_rlt1_i;
    end else begin
      dec_rlt2_o = dec_rlt2_i;
    end
  end

  assign Const_429 = (1'd0 ^ working_key[942]);
  assign Const_430 = (1'd1 ^ working_key[943]);
  assign Const_431 = (1'd1 ^ working_key[944]);

  always @(*) begin
    if(((Const_429 == ap_CS_fsm_state11) ^ working_key[945]) == 1'b1) begin
      dec_rlt2_o_ap_vld = Const_430;
    end else begin
      dec_rlt2_o_ap_vld = Const_431;
    end
  end

  assign Const_432 = (1'd0 ^ working_key[946]);
  assign Const_433 = (1'd1 ^ working_key[947]);

  always @(*) begin
    if(((Const_432 == ap_CS_fsm_state23) ^ working_key[949]) == 1'b0) begin
      grp_upzero_fu_442_bli_q0 = dec_del_bph_q0;
    end else if(((Const_433 == ap_CS_fsm_state12) ^ working_key[948]) == 1'b1) begin
      grp_upzero_fu_442_bli_q0 = dec_del_bpl_q0;
    end else begin
      grp_upzero_fu_442_bli_q0 = 'bx;
    end
  end

  assign Const_434 = (1'd1 ^ working_key[950]);
  assign Const_435 = (1'd0 ^ working_key[951]);

  always @(*) begin
    if(((Const_434 == ap_CS_fsm_state23) ^ working_key[953]) == 1'b0) begin
      grp_upzero_fu_442_dlt = tmp_50_reg_2106;
    end else if(((Const_435 == ap_CS_fsm_state12) ^ working_key[952]) == 1'b1) begin
      grp_upzero_fu_442_dlt = tmp_43_reg_1989;
    end else begin
      grp_upzero_fu_442_dlt = 'bx;
    end
  end

  assign Const_436 = (1'd1 ^ working_key[954]);
  assign Const_437 = (1'd0 ^ working_key[955]);

  always @(*) begin
    if(((Const_436 == ap_CS_fsm_state23) ^ working_key[957]) == 1'b0) begin
      grp_upzero_fu_442_dlti_q0 = dec_del_dhx_q0;
    end else if(((Const_437 == ap_CS_fsm_state12) ^ working_key[956]) == 1'b1) begin
      grp_upzero_fu_442_dlti_q0 = dec_del_dltx_q0;
    end else begin
      grp_upzero_fu_442_dlti_q0 = 'bx;
    end
  end

  assign Const_438 = (1'd1 ^ working_key[958]);
  assign Const_439 = (1'd0 ^ working_key[959]);

  always @(*) begin
    if(((Const_438 == ap_CS_fsm_state23) ^ working_key[961]) == 1'b0) begin
      grp_upzero_fu_442_dlti_q1 = dec_del_dhx_q1;
    end else if(((Const_439 == ap_CS_fsm_state12) ^ working_key[960]) == 1'b1) begin
      grp_upzero_fu_442_dlti_q1 = dec_del_dltx_q1;
    end else begin
      grp_upzero_fu_442_dlti_q1 = 'bx;
    end
  end

  assign Const_440 = (1'd1 ^ working_key[962]);

  always @(*) begin
    if(((Const_440 == ap_CS_fsm_state4) ^ working_key[963]) == 1'b1) begin
      ih_o = ih_i;
    end else begin
      ih_o = ih_assign_fu_529_p1;
    end
  end

  assign Const_441 = (1'd1 ^ working_key[964]);
  assign Const_442 = (1'd0 ^ working_key[965]);
  assign Const_443 = (1'd0 ^ working_key[966]);

  always @(*) begin
    if(((Const_441 == ap_CS_fsm_state4) ^ working_key[967]) == 1'b1) begin
      ih_o_ap_vld = Const_443;
    end else begin
      ih_o_ap_vld = Const_442;
    end
  end

  assign Const_444 = (1'd1 ^ working_key[968]);
  assign Const_445 = (1'd1 ^ working_key[969]);

  always @(*) begin
    if(((Const_444 == ap_CS_fsm_state21) ^ working_key[971]) == 1'b1) begin
      ilb_table_address0 = tmp_i6_fu_1384_p1;
    end else if(((Const_445 == ap_CS_fsm_state10) ^ working_key[970]) == 1'b1) begin
      ilb_table_address0 = tmp_i2_fu_762_p1;
    end else begin
      ilb_table_address0 = 'bx;
    end
  end

  assign Const_446 = (1'd1 ^ working_key[972]);
  assign Const_447 = (1'd0 ^ working_key[973]);
  assign Const_448 = (1'd1 ^ working_key[974]);
  assign Const_449 = (1'd1 ^ working_key[975]);

  always @(*) begin
    if((((Const_446 == ap_CS_fsm_state21) | (Const_447 == ap_CS_fsm_state10)) ^ working_key[976]) == 1'b1) begin
      ilb_table_ce0 = Const_448;
    end else begin
      ilb_table_ce0 = Const_449;
    end
  end

  assign Const_450 = (1'd0 ^ working_key[977]);
  assign Const_451 = (1'd1 ^ working_key[978]);
  assign Const_452 = (1'd1 ^ working_key[979]);

  always @(*) begin
    if(((Const_450 == ap_CS_fsm_state5) ^ working_key[980]) == 1'b1) begin
      qq4_code4_table_ce0 = Const_451;
    end else begin
      qq4_code4_table_ce0 = Const_452;
    end
  end

  assign Const_453 = (1'd0 ^ working_key[981]);
  assign Const_454 = (1'd1 ^ working_key[982]);
  assign Const_455 = (1'd1 ^ working_key[983]);

  always @(*) begin
    if(((Const_453 == ap_CS_fsm_state5) ^ working_key[984]) == 1'b1) begin
      qq6_code6_table_ce0 = Const_454;
    end else begin
      qq6_code6_table_ce0 = Const_455;
    end
  end

  assign Const_456 = (1'd0 ^ working_key[985]);
  assign Const_457 = (1'd1 ^ working_key[986]);
  assign Const_458 = (1'd1 ^ working_key[987]);

  always @(*) begin
    if(((Const_456 == ap_CS_fsm_state5) ^ working_key[988]) == 1'b1) begin
      wl_code_table_ce0 = Const_457;
    end else begin
      wl_code_table_ce0 = Const_458;
    end
  end

  assign Const_459 = (1'd0 ^ working_key[989]);
  assign Const_460 = (1'd1 ^ working_key[990]);
  assign Const_461 = (1'd1 ^ working_key[992]);
  assign Const_462 = (1'd0 ^ working_key[993]);
  assign Const_463 = (1'd1 ^ working_key[995]);
  assign Const_464 = (1'd0 ^ working_key[996]);
  assign Const_465 = (1'd1 ^ working_key[998]);
  assign Const_466 = (1'd1 ^ working_key[999]);
  assign Const_467 = (1'd1 ^ working_key[1001]);
  assign Const_468 = (1'd0 ^ working_key[1002]);
  assign Const_469 = (1'd0 ^ working_key[1004]);
  assign Const_470 = (1'd1 ^ working_key[1005]);

  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if(((ap_start == Const_459) & (Const_460 == ap_CS_fsm_state1) ^ working_key[991]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end
      end
      ap_ST_fsm_state2: begin
        ap_NS_fsm = ap_ST_fsm_state3;
      end
      ap_ST_fsm_state3: begin
        ap_NS_fsm = ap_ST_fsm_state4;
      end
      ap_ST_fsm_state4: begin
        ap_NS_fsm = ap_ST_fsm_state5;
      end
      ap_ST_fsm_state5: begin
        if(((exitcond3_fu_551_p2 == Const_461) & (Const_462 == ap_CS_fsm_state5) ^ working_key[994]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state9;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end
      end
      ap_ST_fsm_state6: begin
        ap_NS_fsm = ap_ST_fsm_state7;
      end
      ap_ST_fsm_state7: begin
        ap_NS_fsm = ap_ST_fsm_state8;
      end
      ap_ST_fsm_state8: begin
        ap_NS_fsm = ap_ST_fsm_state5;
      end
      ap_ST_fsm_state9: begin
        ap_NS_fsm = ap_ST_fsm_state10;
      end
      ap_ST_fsm_state10: begin
        ap_NS_fsm = ap_ST_fsm_state11;
      end
      ap_ST_fsm_state11: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      ap_ST_fsm_state12: begin
        if(((grp_upzero_fu_442_ap_done == Const_463) & (Const_464 == ap_CS_fsm_state12) ^ working_key[997]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state12;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state13;
        end
      end
      ap_ST_fsm_state13: begin
        ap_NS_fsm = ap_ST_fsm_state14;
      end
      ap_ST_fsm_state14: begin
        ap_NS_fsm = ap_ST_fsm_state15;
      end
      ap_ST_fsm_state15: begin
        ap_NS_fsm = ap_ST_fsm_state16;
      end
      ap_ST_fsm_state16: begin
        ap_NS_fsm = ap_ST_fsm_state17;
      end
      ap_ST_fsm_state17: begin
        if(((exitcond2_fu_1202_p2 == Const_465) & (Const_466 == ap_CS_fsm_state17) ^ working_key[1000]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state18;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state21;
        end
      end
      ap_ST_fsm_state18: begin
        ap_NS_fsm = ap_ST_fsm_state19;
      end
      ap_ST_fsm_state19: begin
        ap_NS_fsm = ap_ST_fsm_state20;
      end
      ap_ST_fsm_state20: begin
        ap_NS_fsm = ap_ST_fsm_state17;
      end
      ap_ST_fsm_state21: begin
        ap_NS_fsm = ap_ST_fsm_state22;
      end
      ap_ST_fsm_state22: begin
        ap_NS_fsm = ap_ST_fsm_state23;
      end
      ap_ST_fsm_state23: begin
        if(((grp_upzero_fu_442_ap_done == Const_467) & (Const_468 == ap_CS_fsm_state23) ^ working_key[1003]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state24;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state23;
        end
      end
      ap_ST_fsm_state24: begin
        ap_NS_fsm = ap_ST_fsm_state25;
      end
      ap_ST_fsm_state25: begin
        ap_NS_fsm = ap_ST_fsm_state26;
      end
      ap_ST_fsm_state26: begin
        ap_NS_fsm = ap_ST_fsm_state27;
      end
      ap_ST_fsm_state27: begin
        ap_NS_fsm = ap_ST_fsm_state28;
      end
      ap_ST_fsm_state28: begin
        if(((exitcond_fu_1859_p2 == Const_469) & (Const_470 == ap_CS_fsm_state28) ^ working_key[1006]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state29;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state29: begin
        ap_NS_fsm = ap_ST_fsm_state28;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign ac_ptr_0_sum_cast_fu_1835_p1 = ac_ptr_0_sum_fu_1829_p2;
  assign Const_471 = (5'd31 ^ working_key[1011:1007]);
  assign ac_ptr_0_sum_fu_1829_p2 = (working_key[1012] == 1'b1)? ad_ptr_1_rec_reg_420 << Const_471 : ad_ptr_1_rec_reg_420 + Const_471;
  assign ad_ptr_0_sum7_cast_fu_1853_p1 = ad_ptr_0_sum7_fu_1847_p2;
  assign Const_472 = (5'd27 ^ working_key[1017:1013]);
  assign ad_ptr_0_sum7_fu_1847_p2 = (working_key[1018] == 1'b1)? ad_ptr_1_rec_reg_420 << Const_472 : ad_ptr_1_rec_reg_420 + Const_472;
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];
  assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];
  assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];
  assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];
  assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];
  assign ap_CS_fsm_state21 = ap_CS_fsm[32'd20];
  assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];
  assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];
  assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];
  assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];
  assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];
  assign ap_CS_fsm_state27 = ap_CS_fsm[32'd26];
  assign ap_CS_fsm_state28 = ap_CS_fsm[32'd27];
  assign ap_CS_fsm_state29 = ap_CS_fsm[32'd28];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign apl1_11_cast_fu_1162_p1 = apl1_11_fu_1156_p2;
  assign Const_473 = (16'd23861 ^ working_key[1034:1019]);
  assign apl1_11_fu_1156_p2 = (working_key[1035] == 1'b1)? Const_473 - apl1_17_cast1_fu_1132_p1 : Const_473 << apl1_17_cast1_fu_1132_p1;
  assign apl1_12_cast_fu_1180_p1 = apl1_12_fu_1175_p3;
  assign Const_474 = (1'd1 ^ working_key[1036]);
  assign apl1_12_fu_1175_p3 = ((((working_key[1037] == 1'b1)? tmp_7_i_reg_2047[0:0] === Const_474 : tmp_7_i_reg_2047[0:0] < Const_474) ^ working_key[1038]) == 1'b1)? apl1_11_reg_2042 : tmp_82_reg_2037;
  assign apl1_13_fu_1696_p2 = (working_key[1039] == 1'b1)? tmp7_fu_1690_p2 + tmp_4_i2_cast_cast_fu_1683_p3 : tmp7_fu_1690_p2 >> tmp_4_i2_cast_cast_fu_1683_p3;
  assign apl1_15_cast_fu_1764_p1 = apl1_15_fu_1758_p2;
  assign Const_475 = (16'd21653 ^ working_key[1055:1040]);
  assign apl1_15_fu_1758_p2 = (working_key[1056] == 1'b1)? Const_475 - apl1_18_cast9_fu_1734_p1 : Const_475 + apl1_18_cast9_fu_1734_p1;
  assign apl1_16_cast_fu_1784_p1 = apl1_16_fu_1779_p3;
  assign Const_476 = (1'd0 ^ working_key[1057]);
  assign apl1_16_fu_1779_p3 = ((((working_key[1058] == 1'b1)? tmp_7_i2_reg_2186[0:0] == Const_476 : tmp_7_i2_reg_2186[0:0] === Const_476) ^ working_key[1059]) == 1'b1)? apl1_15_reg_2181 : tmp_95_reg_2176;
  assign apl1_17_cast1_fu_1132_p1 = apl1_17_fu_1127_p2;
  assign apl1_17_cast_fu_1136_p1 = apl1_17_fu_1127_p2;
  assign Const_477 = (15'd27133 ^ working_key[1074:1060]);
  assign apl1_17_fu_1127_p2 = (working_key[1075] == 1'b1)? Const_477 * apl2_assign_reg_2025 : Const_477 - apl2_assign_reg_2025;
  assign apl1_18_cast9_fu_1734_p1 = apl1_18_fu_1729_p2;
  assign apl1_18_cast_fu_1738_p1 = apl1_18_fu_1729_p2;
  assign Const_478 = (15'd5802 ^ working_key[1090:1076]);
  assign apl1_18_fu_1729_p2 = (working_key[1091] == 1'b1)? Const_478 - apl2_assign_2_reg_2164 : Const_478 << apl2_assign_2_reg_2164;
  assign apl1_fu_1112_p2 = (working_key[1092] == 1'b1)? tmp_4_i_cast_cast_fu_1099_p3 - tmp5_fu_1106_p2 : tmp_4_i_cast_cast_fu_1099_p3 + tmp5_fu_1106_p2;
  assign apl2_2_fu_1606_p2 = (working_key[1093] == 1'b1)? tmp6_cast_fu_1602_p1 + tmp_8_i2_cast_cast_fu_1562_p3 : tmp6_cast_fu_1602_p1 - tmp_8_i2_cast_cast_fu_1562_p3;
  assign apl2_assign_2_cast_fu_1720_p1 = apl2_assign_2_reg_2164;
  assign Const_479 = (1'd1 ^ working_key[1094]);
  assign Const_480 = (15'd31392 ^ working_key[1110:1096]);
  assign apl2_assign_2_fu_1672_p3 = ((((working_key[1095] == 1'b1)? tmp_3_i2_fu_1666_p2[0:0] === Const_479 : tmp_3_i2_fu_1666_p2[0:0] != Const_479) ^ working_key[1111]) == 1'b1)? tmp_92_fu_1662_p1 : Const_480;
  assign apl2_assign_cast_fu_1118_p1 = apl2_assign_reg_2025;
  assign Const_481 = (1'd1 ^ working_key[1112]);
  assign Const_482 = (15'd15530 ^ working_key[1128:1114]);
  assign apl2_assign_fu_1088_p3 = ((((working_key[1113] == 1'b1)? tmp_3_i_fu_1082_p2[0:0] === Const_481 : tmp_3_i_fu_1082_p2[0:0] != Const_481) ^ working_key[1129]) == 1'b1)? tmp_79_fu_1078_p1 : Const_482;
  assign apl2_fu_1038_p2 = (working_key[1130] == 1'b1)? tmp_8_i_cast_cast_fu_994_p3 + tmp4_cast_fu_1034_p1 : tmp_8_i_cast_cast_fu_994_p3 << tmp4_cast_fu_1034_p1;
  assign dec_del_bph_d0 = grp_upzero_fu_442_bli_d0;
  assign dec_del_bpl_d0 = grp_upzero_fu_442_bli_d0;
  assign dec_del_dhx_address1 = grp_upzero_fu_442_dlti_address1;
  assign dec_del_dhx_d0 = grp_upzero_fu_442_dlti_d0;
  assign dec_del_dhx_d1 = grp_upzero_fu_442_dlti_d1;
  assign dec_del_dltx_address1 = grp_upzero_fu_442_dlti_address1;
  assign dec_del_dltx_d0 = grp_upzero_fu_442_dlti_d0;
  assign dec_del_dltx_d1 = grp_upzero_fu_442_dlti_d1;
  assign dec_rlt_fu_874_p2 = (working_key[1131] == 1'b1)? dec_sl_cast_fu_805_p1 * dec_dlt : dec_sl_cast_fu_805_p1 + dec_dlt;
  assign dec_sl_cast_fu_805_p1 = dec_sl_fu_799_p2;
  assign dec_sl_fu_799_p2 = (working_key[1132] == 1'b1)? tmp_20_i_cast_fu_795_p1 + tmp_i_cast_fu_777_p1 : tmp_20_i_cast_fu_795_p1 * tmp_i_cast_fu_777_p1;
  assign dl_cast_fu_816_p1 = tmp_71_reg_1974;
  assign Const_483 = (3'd3 ^ working_key[1135:1133]);
  assign Const_484 = (1'd0 ^ working_key[1137]);
  assign Const_485 = (1'd0 ^ working_key[1138]);
  assign exitcond2_fu_1202_p2 = ((((working_key[1136] == 1'b1)? dlt_pn_rec_i2_reg_409 > Const_483 : dlt_pn_rec_i2_reg_409 == Const_483) ^ working_key[1139]) == 1'b1)? Const_485 : Const_484;
  assign Const_486 = (3'd1 ^ working_key[1142:1140]);
  assign Const_487 = (1'd1 ^ working_key[1144]);
  assign Const_488 = (1'd1 ^ working_key[1145]);
  assign exitcond3_fu_551_p2 = ((((working_key[1143] == 1'b1)? dlt_pn_rec_i_reg_388 === Const_486 : dlt_pn_rec_i_reg_388 == Const_486) ^ working_key[1146]) == 1'b1)? Const_487 : Const_488;
  assign Const_489 = (4'd15 ^ working_key[1150:1147]);
  assign Const_490 = (1'd0 ^ working_key[1152]);
  assign Const_491 = (1'd0 ^ working_key[1153]);
  assign exitcond_fu_1859_p2 = ((((working_key[1151] == 1'b1)? i_1_reg_431 == Const_489 : i_1_reg_431 > Const_489) ^ working_key[1154]) == 1'b1)? Const_490 : Const_491;
  assign extLd_cast_fu_670_p1 = dec_detl_i;
  assign grp_fu_493_p2 = (working_key[1155] == 1'b1)? reg_489 * reg_485 : reg_489 << reg_485;
  assign grp_upzero_fu_442_ap_start = grp_upzero_fu_442_ap_start_reg;
  assign Const_492 = (4'd15 ^ working_key[1159:1156]);
  assign i_fu_1865_p2 = (working_key[1160] == 1'b1)? i_1_reg_431 - Const_492 : i_1_reg_431 + Const_492;
  assign ih_assign_fu_529_p1 = tmp_41_fu_519_p4;
  assign nbh_assign_2_cast_fu_1288_p2 = (working_key[1161] == 1'b1)? tmp_16_fu_1274_p1 + tmp_85_fu_1278_p1 : tmp_16_fu_1274_p1 - tmp_85_fu_1278_p1;
  assign nbh_assign_2_fu_1282_p2 = (working_key[1162] == 1'b1)? tmp_15_fu_1260_p6 * wd_fu_1256_p1 : tmp_15_fu_1260_p6 + wd_fu_1256_p1;
  assign nbl_assign_4_cast_fu_636_p2 = (working_key[1163] == 1'b1)? tmp_13_fu_626_p1 + tmp_32_i_fu_608_p4 : tmp_13_fu_626_p1 * tmp_32_i_fu_608_p4;
  assign nbl_assign_4_fu_630_p2 = (working_key[1164] == 1'b1)? wd_cast_fu_618_p1 - wl_code_table_load_c_fu_622_p1 : wd_cast_fu_618_p1 + wl_code_table_load_c_fu_622_p1;
  assign nbl_assign_5_cast_fu_732_p1 = nbl_assign_5_fu_724_p3;
  assign Const_493 = (1'd0 ^ working_key[1165]);
  assign Const_494 = (15'd24875 ^ working_key[1181:1167]);
  assign nbl_assign_5_fu_724_p3 = ((((working_key[1166] == 1'b1)? tmp_18_i_fu_718_p2[0:0] == Const_493 : tmp_18_i_fu_718_p2[0:0] === Const_493) ^ working_key[1182]) == 1'b1)? tmp_74_fu_714_p1 : Const_494;
  assign nbl_assign_6_cast_fu_1354_p1 = nbl_assign_6_fu_1346_p3;
  assign Const_495 = (1'd1 ^ working_key[1183]);
  assign Const_496 = (15'd30697 ^ working_key[1199:1185]);
  assign nbl_assign_6_fu_1346_p3 = ((((working_key[1184] == 1'b1)? tmp_19_i3_fu_1340_p2[0:0] === Const_495 : tmp_19_i3_fu_1340_p2[0:0] == Const_495) ^ working_key[1200]) == 1'b1)? tmp_87_fu_1336_p1 : Const_496;
  assign p_01_rec_i2_cast_fu_1196_p1 = p_01_rec_i2_fu_1190_p2;
  assign Const_497 = (3'd3 ^ working_key[1203:1201]);
  assign p_01_rec_i2_fu_1190_p2 = (working_key[1204] == 1'b1)? dlt_pn_rec_i2_reg_409 << Const_497 : dlt_pn_rec_i2_reg_409 + Const_497;
  assign p_01_rec_i_cast_fu_545_p1 = p_01_rec_i_fu_539_p2;
  assign Const_498 = (3'd4 ^ working_key[1207:1205]);
  assign p_01_rec_i_fu_539_p2 = (working_key[1208] == 1'b1)? dlt_pn_rec_i_reg_388 >> Const_498 : dlt_pn_rec_i_reg_388 + Const_498;
  assign Const_499 = (1'd0 ^ working_key[1209]);
  assign Const_500 = (27'd89400661 ^ working_key[1237:1211]);
  assign p_i4_fu_1071_p3 = ((((working_key[1210] == 1'b1)? tmp_2_i_fu_1066_p2[0:0] < Const_499 : tmp_2_i_fu_1066_p2[0:0] === Const_499) ^ working_key[1238]) == 1'b1)? Const_500 : apl2_reg_2014;
  assign Const_501 = (1'd0 ^ working_key[1239]);
  assign Const_502 = (31'd627743061 ^ working_key[1271:1241]);
  assign p_i5_fu_1330_p3 = ((((working_key[1240] == 1'b1)? tmp_86_reg_2091[0:0] > Const_501 : tmp_86_reg_2091[0:0] === Const_501) ^ working_key[1272]) == 1'b1)? Const_502 : nbh_assign_2_cast_reg_2086;
  assign Const_503 = (1'd0 ^ working_key[1273]);
  assign Const_504 = (27'd45444405 ^ working_key[1301:1275]);
  assign p_i6_fu_1655_p3 = ((((working_key[1274] == 1'b1)? tmp_2_i2_fu_1650_p2[0:0] == Const_503 : tmp_2_i2_fu_1650_p2[0:0] === Const_503) ^ working_key[1302]) == 1'b1)? Const_504 : apl2_2_reg_2143;
  assign Const_505 = (1'd0 ^ working_key[1303]);
  assign Const_506 = (25'd11528618 ^ working_key[1329:1305]);
  assign p_i_fu_708_p3 = ((((working_key[1304] == 1'b1)? tmp_73_reg_1953[0:0] != Const_505 : tmp_73_reg_1953[0:0] === Const_505) ^ working_key[1330]) == 1'b1)? nbl_assign_4_cast_reg_1948 : Const_506;
  assign Const_507 = (5'd11 ^ working_key[1335:1331]);
  assign p_rec_fu_1841_p2 = (working_key[1336] == 1'b1)? ad_ptr_1_rec_reg_420 << Const_507 : ad_ptr_1_rec_reg_420 + Const_507;
  assign pl_2_fu_1638_p0 = dec_ah1_i;
  assign pl_2_fu_1638_p1 = dec_rh1_i;
  assign pl_2_fu_1638_p2 = (working_key[1337] == 1'b1)? pl_2_fu_1638_p0 * pl_2_fu_1638_p1 : pl_2_fu_1638_p0 - pl_2_fu_1638_p1;
  assign pl_fu_654_p0 = dec_rlt1_i;
  assign pl_fu_654_p1 = dec_al1_i;
  assign pl_fu_654_p2 = (working_key[1338] == 1'b1)? pl_fu_654_p0 << pl_fu_654_p1 : pl_fu_654_p0 * pl_fu_654_p1;
  assign qq4_code4_table_address0 = tmp_s_fu_566_p1;
  assign qq6_code6_table_address0 = tmp_45_fu_576_p1;
  assign rh_fu_1801_p2 = (working_key[1339] == 1'b1)? tmp8_cast_fu_1798_p1 + dec_dh : tmp8_cast_fu_1798_p1 >> dec_dh;
  assign rl_cast_fu_1172_p1 = rl_reg_1994;
  assign rl_fu_819_p2 = (working_key[1340] == 1'b1)? dl_cast_fu_816_p1 * dec_sl_fu_799_p2 : dl_cast_fu_816_p1 + dec_sl_fu_799_p2;
  assign tmp4_cast_fu_1034_p1 = tmp4_fu_1028_p2;
  assign tmp4_fu_1028_p2 = (working_key[1341] == 1'b1)? wd2_15_cast_fu_983_p1 + tmp_1_i_cast_fu_1024_p1 : wd2_15_cast_fu_983_p1 * tmp_1_i_cast_fu_1024_p1;
  assign Const_508 = (25'd11174506 ^ working_key[1366:1342]);
  assign tmp5_fu_1106_p2 = (working_key[1367] == 1'b1)? Const_508 + wd2_16_cast_fu_1096_p1 : Const_508 >> wd2_16_cast_fu_1096_p1;
  assign tmp6_cast_fu_1602_p1 = tmp6_fu_1596_p2;
  assign tmp6_fu_1596_p2 = (working_key[1368] == 1'b1)? tmp_1_i2_cast_fu_1592_p1 - wd2_21_cast_fu_1551_p1 : tmp_1_i2_cast_fu_1592_p1 + wd2_21_cast_fu_1551_p1;
  assign Const_509 = (25'd5675413 ^ working_key[1393:1369]);
  assign tmp7_fu_1690_p2 = (working_key[1394] == 1'b1)? Const_509 + wd2_22_cast_fu_1680_p1 : Const_509 * wd2_22_cast_fu_1680_p1;
  assign tmp8_cast_fu_1798_p1 = tmp8_reg_2191;
  assign tmp8_fu_1774_p2 = (working_key[1395] == 1'b1)? tmp_i19_cast_reg_2123 << tmp_20_i5_cast_fu_1716_p1 : tmp_i19_cast_reg_2123 + tmp_20_i5_cast_fu_1716_p1;
  assign tmp_10_i2_fu_1430_p3 = { { wd3_5_fu_1424_p2 }, { 3'd0 } };
  assign tmp_10_i_fu_840_p3 = { { wd3_fu_834_p2 }, { 3'd0 } };
  assign tmp_13_fu_626_p0 = wl_code_table_q0;
  assign tmp_13_fu_626_p1 = tmp_13_fu_626_p0;
  assign tmp_16_fu_1274_p1 = tmp_36_i_fu_1246_p4;
  assign Const_510 = (25'd27959722 ^ working_key[1420:1396]);
  assign Const_511 = (1'd0 ^ working_key[1422]);
  assign Const_512 = (1'd0 ^ working_key[1423]);
  assign tmp_18_i_fu_718_p2 = ((((working_key[1421] == 1'b1)? p_i_fu_708_p3 < Const_510 : p_i_fu_708_p3 > Const_510) ^ working_key[1424]) == 1'b1)? Const_512 : Const_511;
  assign Const_513 = (31'd721339044 ^ working_key[1455:1425]);
  assign Const_514 = (1'd0 ^ working_key[1457]);
  assign Const_515 = (1'd0 ^ working_key[1458]);
  assign tmp_19_i3_fu_1340_p2 = ((((working_key[1456] == 1'b1)? p_i5_fu_1330_p3 < Const_513 : p_i5_fu_1330_p3 > Const_513) ^ working_key[1459]) == 1'b1)? Const_515 : Const_514;
  assign tmp_19_i4_fu_1582_p4 = { { tmp_9_i6_fu_1576_p2[31:7] } };
  assign tmp_19_i_fu_1014_p4 = { { tmp_9_i4_fu_1008_p2[31:7] } };
  assign tmp_1_cast_fu_557_p4 = { { input_r[5:2] } };
  assign tmp_1_i2_cast_fu_1592_p1 = tmp_19_i4_fu_1582_p4;
  assign tmp_1_i_cast_fu_1024_p1 = tmp_19_i_fu_1014_p4;
  assign tmp_20_i5_cast_fu_1716_p1 = tmp_41_i2_fu_1706_p4;
  assign tmp_20_i_cast_fu_795_p1 = tmp_41_i_fu_785_p4;
  assign Const_516 = (27'd44079786 ^ working_key[1486:1460]);
  assign Const_517 = (1'd1 ^ working_key[1488]);
  assign Const_518 = (1'd1 ^ working_key[1489]);
  assign tmp_2_i2_fu_1650_p2 = ((((working_key[1487] == 1'b1)? apl2_2_reg_2143 > Const_516 : apl2_2_reg_2143 < Const_516) ^ working_key[1490]) == 1'b1)? Const_517 : Const_518;
  assign Const_519 = (27'd95049045 ^ working_key[1517:1491]);
  assign Const_520 = (1'd0 ^ working_key[1519]);
  assign Const_521 = (1'd0 ^ working_key[1520]);
  assign tmp_2_i_fu_1066_p2 = ((((working_key[1518] == 1'b1)? apl2_reg_2014 != Const_519 : apl2_reg_2014 > Const_519) ^ working_key[1521]) == 1'b1)? Const_520 : Const_521;
  assign tmp_32_i_fu_608_p4 = { { tmp_i7_fu_602_p2[31:7] } };
  assign tmp_36_i_fu_1246_p4 = { { tmp_i2_35_fu_1240_p2[31:7] } };
  assign tmp_39_i2_fu_1389_p4 = { { zl1_i2_reg_399[31:14] } };
  assign tmp_39_i_fu_767_p4 = { { zl1_i_reg_378[31:14] } };
  assign Const_522 = (27'd22312617 ^ working_key[1548:1522]);
  assign Const_523 = (1'd0 ^ working_key[1550]);
  assign Const_524 = (1'd0 ^ working_key[1551]);
  assign tmp_3_i2_fu_1666_p2 = ((((working_key[1549] == 1'b1)? p_i6_fu_1655_p3 > Const_522 : p_i6_fu_1655_p3 < Const_522) ^ working_key[1552]) == 1'b1)? Const_524 : Const_523;
  assign Const_525 = (27'd83970724 ^ working_key[1579:1553]);
  assign Const_526 = (1'd1 ^ working_key[1581]);
  assign Const_527 = (1'd1 ^ working_key[1582]);
  assign tmp_3_i_fu_1082_p2 = ((((working_key[1580] == 1'b1)? p_i4_fu_1071_p3 < Const_525 : p_i4_fu_1071_p3 == Const_525) ^ working_key[1583]) == 1'b1)? Const_526 : Const_527;
  assign tmp_41_fu_519_p4 = { { input_r[31:6] } };
  assign tmp_41_i2_fu_1706_p4 = { { tmp_i1_34_fu_1702_p2[30:14] } };
  assign tmp_41_i_fu_785_p4 = { { tmp_i_31_fu_781_p2[30:14] } };
  assign tmp_42_fu_1871_p1 = extLd_cast_fu_670_p1;
  assign tmp_43_fu_809_p1 = tmp_70_reg_1968;
  assign tmp_44_fu_686_p1 = tmp_70_fu_677_p4;
  assign tmp_45_fu_576_p1 = il;
  assign tmp_46_fu_1878_p1 = extLd_cast_fu_670_p1;
  assign tmp_48_fu_854_p2 = (working_key[1584] == 1'b1)? tmp_59_cast_fu_813_p1 >> tmp_i_cast_fu_777_p1 : tmp_59_cast_fu_813_p1 + tmp_i_cast_fu_777_p1;
  assign tmp_49_fu_1315_p0 = tmp_49_fu_1315_p00;
  assign tmp_49_fu_1315_p00 = dec_deth_i;
  assign Const_528 = (32'd1426412885 ^ working_key[1616:1585]);
  assign tmp_49_fu_1315_p2 = (working_key[1617] == 1'b1)? { { Const_528 }, { tmp_49_fu_1315_p0 } } * tmp_14_reg_2081 : { { Const_528 }, { tmp_49_fu_1315_p0 } } - tmp_14_reg_2081;
  assign Const_529 = (1'd1 ^ working_key[1618]);
  assign Const_530 = (25'd19418154 ^ working_key[1644:1620]);
  assign Const_531 = (25'd24433957 ^ working_key[1669:1645]);
  assign tmp_4_i2_cast_cast_fu_1683_p3 = ((((working_key[1619] == 1'b1)? tmp_94_reg_2138[0:0] === Const_529 : tmp_94_reg_2138[0:0] > Const_529) ^ working_key[1670]) == 1'b1)? Const_530 : Const_531;
  assign Const_532 = (1'd0 ^ working_key[1671]);
  assign Const_533 = (25'd23419437 ^ working_key[1697:1673]);
  assign Const_534 = (25'd11179391 ^ working_key[1722:1698]);
  assign tmp_4_i_cast_cast_fu_1099_p3 = ((((working_key[1672] == 1'b1)? tmp_81_reg_2009[0:0] > Const_532 : tmp_81_reg_2009[0:0] === Const_532) ^ working_key[1723]) == 1'b1)? Const_534 : Const_533;
  assign tmp_51_fu_1403_p1 = tmp_50_reg_2106;
  assign tmp_52_fu_1444_p2 = (working_key[1724] == 1'b1)? tmp_i19_cast_fu_1399_p1 - tmp_69_cast_fu_1406_p1 : tmp_i19_cast_fu_1399_p1 + tmp_69_cast_fu_1406_p1;
  assign tmp_53_fu_955_p4 = { { wd2_4_fu_949_p2[31:7] } };
  assign tmp_54_fu_965_p4 = { { dec_al1_i[29:5] } };
  assign Const_535 = (1'd0 ^ working_key[1725]);
  assign tmp_55_fu_975_p3 = ((((working_key[1726] == 1'b1)? tmp_76_fu_942_p3[0:0] < Const_535 : tmp_76_fu_942_p3[0:0] === Const_535) ^ working_key[1727]) == 1'b1)? tmp_53_fu_955_p4 : tmp_54_fu_965_p4;
  assign tmp_56_fu_1523_p4 = { { wd2_6_fu_1517_p2[31:7] } };
  assign tmp_57_fu_1533_p4 = { { dec_ah1_i[29:5] } };
  assign Const_536 = (1'd1 ^ working_key[1728]);
  assign tmp_58_fu_1543_p3 = ((((working_key[1729] == 1'b1)? tmp_89_fu_1510_p3[0:0] === Const_536 : tmp_89_fu_1510_p3[0:0] == Const_536) ^ working_key[1730]) == 1'b1)? tmp_57_fu_1533_p4 : tmp_56_fu_1523_p4;
  assign tmp_59_cast_fu_813_p1 = tmp_70_reg_1968;
  assign tmp_5_i5_fu_1478_p0 = dec_ph;
  assign tmp_5_i5_fu_1478_p1 = dec_ph2_i;
  assign tmp_5_i5_fu_1478_p2 = (working_key[1731] == 1'b1)? tmp_5_i5_fu_1478_p0 * tmp_5_i5_fu_1478_p1 : tmp_5_i5_fu_1478_p0 + tmp_5_i5_fu_1478_p1;
  assign tmp_5_i_fu_910_p0 = dec_plt2_i;
  assign tmp_5_i_fu_910_p1 = dec_plt;
  assign tmp_5_i_fu_910_p2 = (working_key[1732] == 1'b1)? tmp_5_i_fu_910_p0 >> tmp_5_i_fu_910_p1 : tmp_5_i_fu_910_p0 * tmp_5_i_fu_910_p1;
  assign tmp_64_cast_fu_860_p1 = tmp_48_fu_854_p2;
  assign tmp_69_cast_fu_1406_p1 = tmp_50_reg_2106;
  assign Const_537 = (1'd1 ^ working_key[1734]);
  assign Const_538 = (1'd0 ^ working_key[1735]);
  assign tmp_6_i2_fu_1742_p2 = ((((working_key[1733] == 1'b1)? apl1_13_reg_2170 < apl1_18_cast_fu_1738_p1 : apl1_13_reg_2170 > apl1_18_cast_fu_1738_p1) ^ working_key[1736]) == 1'b1)? Const_537 : Const_538;
  assign Const_539 = (1'd1 ^ working_key[1738]);
  assign Const_540 = (1'd1 ^ working_key[1739]);
  assign tmp_6_i_fu_1140_p2 = ((((working_key[1737] == 1'b1)? apl1_reg_2031 > apl1_17_cast_fu_1136_p1 : apl1_reg_2031 != apl1_17_cast_fu_1136_p1) ^ working_key[1740]) == 1'b1)? Const_539 : Const_540;
  assign tmp_70_cast_fu_1450_p1 = tmp_52_fu_1444_p2;
  assign tmp_70_fu_677_p4 = { { tmp_42_fu_1871_p2[30:15] } };
  assign Const_541 = (32'd1788433746 ^ working_key[1772:1741]);
  assign tmp_72_fu_596_p2 = (working_key[1773] == 1'b1)? dec_nbl_i << Const_541 : dec_nbl_i >> Const_541;
  assign tmp_74_fu_714_p1 = p_i_fu_708_p3[14:0];
  assign tmp_76_fu_942_p3 = tmp_i8_reg_1999[32'd31];
  assign tmp_77_fu_987_p3 = tmp_5_i_reg_2004[32'd31];
  assign Const_542 = (32'd1790601877 ^ working_key[1805:1774]);
  assign tmp_78_fu_1002_p2 = (working_key[1806] == 1'b1)? dec_al2_i << Const_542 : dec_al2_i >> Const_542;
  assign tmp_79_fu_1078_p1 = p_i4_fu_1071_p3[14:0];
  assign Const_543 = (1'd0 ^ working_key[1808]);
  assign Const_544 = (1'd0 ^ working_key[1809]);
  assign tmp_7_i2_fu_1768_p2 = ((((working_key[1807] == 1'b1)? wd3_0_apl1_i2_fu_1747_p3 > apl1_15_cast_fu_1764_p1 : wd3_0_apl1_i2_fu_1747_p3 < apl1_15_cast_fu_1764_p1) ^ working_key[1810]) == 1'b1)? Const_543 : Const_544;
  assign Const_545 = (1'd1 ^ working_key[1812]);
  assign Const_546 = (1'd0 ^ working_key[1813]);
  assign tmp_7_i_fu_1166_p2 = ((((working_key[1811] == 1'b1)? wd3_0_apl1_i_fu_1145_p3 < apl1_11_cast_fu_1162_p1 : wd3_0_apl1_i_fu_1145_p3 === apl1_11_cast_fu_1162_p1) ^ working_key[1814]) == 1'b1)? Const_546 : Const_545;
  assign Const_547 = (32'd1420556898 ^ working_key[1846:1815]);
  assign tmp_80_fu_1044_p2 = (working_key[1847] == 1'b1)? dec_al1_i << Const_547 : dec_al1_i >> Const_547;
  assign tmp_82_fu_1152_p1 = wd3_0_apl1_i_fu_1145_p3[15:0];
  assign tmp_83_fu_1212_p1 = ih_i[1:0];
  assign Const_548 = (32'd2863270573 ^ working_key[1879:1848]);
  assign tmp_84_fu_1234_p2 = (working_key[1880] == 1'b1)? dec_nbh_i >> Const_548 : dec_nbh_i << Const_548;
  assign tmp_85_fu_1278_p1 = tmp_15_fu_1260_p6[30:0];
  assign tmp_87_fu_1336_p1 = p_i5_fu_1330_p3[14:0];
  assign tmp_89_fu_1510_p3 = tmp_i3_reg_2128[32'd31];
  assign Const_549 = (1'd0 ^ working_key[1881]);
  assign Const_550 = (27'd57299173 ^ working_key[1909:1883]);
  assign Const_551 = (27'd90880746 ^ working_key[1936:1910]);
  assign tmp_8_i2_cast_cast_fu_1562_p3 = ((((working_key[1882] == 1'b1)? tmp_90_fu_1555_p3[0:0] == Const_549 : tmp_90_fu_1555_p3[0:0] === Const_549) ^ working_key[1937]) == 1'b1)? Const_550 : Const_551;
  assign Const_552 = (1'd1 ^ working_key[1938]);
  assign Const_553 = (27'd44051668 ^ working_key[1966:1940]);
  assign Const_554 = (27'd68507092 ^ working_key[1993:1967]);
  assign tmp_8_i_cast_cast_fu_994_p3 = ((((working_key[1939] == 1'b1)? tmp_77_fu_987_p3[0:0] === Const_552 : tmp_77_fu_987_p3[0:0] != Const_552) ^ working_key[1994]) == 1'b1)? Const_553 : Const_554;
  assign tmp_90_fu_1555_p3 = tmp_5_i5_reg_2133[32'd31];
  assign Const_555 = (32'd2858767698 ^ working_key[2026:1995]);
  assign tmp_91_fu_1570_p2 = (working_key[2027] == 1'b1)? dec_ah2_i << Const_555 : dec_ah2_i >> Const_555;
  assign tmp_92_fu_1662_p1 = p_i6_fu_1655_p3[14:0];
  assign Const_556 = (32'd2867440194 ^ working_key[2059:2028]);
  assign tmp_93_fu_1612_p2 = (working_key[2060] == 1'b1)? dec_ah1_i << Const_556 : dec_ah1_i >> Const_556;
  assign tmp_95_fu_1754_p1 = wd3_0_apl1_i2_fu_1747_p3[15:0];
  assign tmp_9_i4_fu_1008_p2 = (working_key[2061] == 1'b1)? tmp_78_fu_1002_p2 >> dec_al2_i : tmp_78_fu_1002_p2 - dec_al2_i;
  assign tmp_9_i5_cast_cast_fu_1420_p1 = tmp_9_i5_fu_1415_p2;
  assign Const_557 = (4'd14 ^ working_key[2065:2062]);
  assign tmp_9_i5_fu_1415_p2 = (working_key[2066] == 1'b1)? Const_557 + wd2_17_cast_reg_2113 : Const_557 - wd2_17_cast_reg_2113;
  assign tmp_9_i6_fu_1576_p2 = (working_key[2067] == 1'b1)? tmp_91_fu_1570_p2 - dec_ah2_i : tmp_91_fu_1570_p2 >> dec_ah2_i;
  assign tmp_9_i_cast_cast_fu_830_p1 = tmp_9_i_fu_825_p2;
  assign Const_558 = (4'd13 ^ working_key[2071:2068]);
  assign tmp_9_i_fu_825_p2 = (working_key[2072] == 1'b1)? Const_558 - wd2_cast_reg_1979 : Const_558 + wd2_cast_reg_1979;
  assign tmp_i19_cast_fu_1399_p1 = tmp_39_i2_fu_1389_p4;
  assign tmp_i1_34_fu_1702_p2 = (working_key[2073] == 1'b1)? tmp_i4_reg_2159 - pl_2_reg_2154 : tmp_i4_reg_2159 + pl_2_reg_2154;
  assign tmp_i1_fu_660_p0 = dec_rlt2_i;
  assign tmp_i1_fu_660_p1 = dec_al2_i;
  assign tmp_i1_fu_660_p2 = (working_key[2074] == 1'b1)? tmp_i1_fu_660_p0 * tmp_i1_fu_660_p1 : tmp_i1_fu_660_p0 + tmp_i1_fu_660_p1;
  assign tmp_i2_35_fu_1240_p2 = (working_key[2075] == 1'b1)? tmp_84_fu_1234_p2 * dec_nbh_i : tmp_84_fu_1234_p2 - dec_nbh_i;
  assign tmp_i2_fu_762_p1 = wd1_fu_742_p4;
  assign tmp_i3_fu_1472_p0 = dec_ph;
  assign tmp_i3_fu_1472_p1 = dec_ph1_i;
  assign tmp_i3_fu_1472_p2 = (working_key[2076] == 1'b1)? tmp_i3_fu_1472_p0 * tmp_i3_fu_1472_p1 : tmp_i3_fu_1472_p0 >> tmp_i3_fu_1472_p1;
  assign tmp_i4_36_fu_1618_p2 = (working_key[2077] == 1'b1)? tmp_93_fu_1612_p2 - dec_ah1_i : tmp_93_fu_1612_p2 * dec_ah1_i;
  assign tmp_i4_fu_1644_p0 = dec_ah2_i;
  assign tmp_i4_fu_1644_p1 = dec_rh2_i;
  assign tmp_i4_fu_1644_p2 = (working_key[2078] == 1'b1)? tmp_i4_fu_1644_p0 << tmp_i4_fu_1644_p1 : tmp_i4_fu_1644_p0 * tmp_i4_fu_1644_p1;
  assign tmp_i6_fu_1384_p1 = wd1_2_fu_1364_p4;
  assign tmp_i7_fu_602_p2 = (working_key[2079] == 1'b1)? tmp_72_fu_596_p2 >> dec_nbl_i : tmp_72_fu_596_p2 - dec_nbl_i;
  assign tmp_i8_fu_904_p0 = dec_plt1_i;
  assign tmp_i8_fu_904_p1 = dec_plt;
  assign tmp_i8_fu_904_p2 = (working_key[2080] == 1'b1)? tmp_i8_fu_904_p0 * tmp_i8_fu_904_p1 : tmp_i8_fu_904_p0 << tmp_i8_fu_904_p1;
  assign tmp_i9_fu_1050_p2 = (working_key[2081] == 1'b1)? tmp_80_fu_1044_p2 + dec_al1_i : tmp_80_fu_1044_p2 - dec_al1_i;
  assign tmp_i_31_fu_781_p2 = (working_key[2082] == 1'b1)? pl_reg_1958 + tmp_i1_reg_1963 : pl_reg_1958 - tmp_i1_reg_1963;
  assign tmp_i_cast_fu_777_p1 = tmp_39_i_fu_767_p4;
  assign tmp_i_fu_581_p2 = (working_key[2083] == 1'b1)? reg_481 * reg_477 : reg_481 + reg_477;
  assign tmp_s_fu_566_p1 = tmp_1_cast_fu_557_p4;
  assign wd1_2_fu_1364_p4 = { { nbl_assign_6_fu_1346_p3[10:6] } };
  assign wd1_fu_742_p4 = { { nbl_assign_5_fu_724_p3[10:6] } };
  assign wd2_15_cast_fu_983_p1 = tmp_55_fu_975_p3;
  assign wd2_16_cast_fu_1096_p1 = tmp_21_i_reg_2020;
  assign wd2_21_cast_fu_1551_p1 = tmp_58_fu_1543_p3;
  assign wd2_22_cast_fu_1680_p1 = tmp_21_i2_reg_2149;
  assign Const_559 = (32'd2863310175 ^ working_key[2115:2084]);
  assign wd2_4_fu_949_p2 = (working_key[2116] == 1'b1)? Const_559 + wd2_fu_936_p2 : Const_559 - wd2_fu_936_p2;
  assign Const_560 = (32'd3646248274 ^ working_key[2148:2117]);
  assign wd2_5_fu_1504_p2 = (working_key[2149] == 1'b1)? dec_ah1_i << Const_560 : dec_ah1_i >> Const_560;
  assign Const_561 = (32'd3127546549 ^ working_key[2181:2150]);
  assign wd2_6_fu_1517_p2 = (working_key[2182] == 1'b1)? Const_561 << wd2_5_fu_1504_p2 : Const_561 - wd2_5_fu_1504_p2;
  assign Const_562 = (32'd4201288375 ^ working_key[2214:2183]);
  assign wd2_fu_936_p2 = (working_key[2215] == 1'b1)? dec_al1_i << Const_562 : dec_al1_i >> Const_562;
  assign Const_563 = (1'd0 ^ working_key[2216]);
  assign wd3_0_apl1_i2_fu_1747_p3 = ((((working_key[2217] == 1'b1)? tmp_6_i2_fu_1742_p2[0:0] != Const_563 : tmp_6_i2_fu_1742_p2[0:0] === Const_563) ^ working_key[2218]) == 1'b1)? apl1_13_reg_2170 : apl1_18_cast_fu_1738_p1;
  assign Const_564 = (1'd1 ^ working_key[2219]);
  assign wd3_0_apl1_i_fu_1145_p3 = ((((working_key[2220] == 1'b1)? tmp_6_i_fu_1140_p2[0:0] === Const_564 : tmp_6_i_fu_1140_p2[0:0] == Const_564) ^ working_key[2221]) == 1'b1)? apl1_17_cast_fu_1136_p1 : apl1_reg_2031;
  assign wd3_5_fu_1424_p2 = (working_key[2222] == 1'b1)? ilb_table_q0 >> tmp_9_i5_cast_cast_fu_1420_p1 : ilb_table_q0 << tmp_9_i5_cast_cast_fu_1420_p1;
  assign wd3_fu_834_p2 = (working_key[2223] == 1'b1)? ilb_table_q0 << tmp_9_i_cast_cast_fu_830_p1 : ilb_table_q0 >> tmp_9_i_cast_cast_fu_830_p1;
  assign wd_cast_fu_618_p1 = tmp_32_i_fu_608_p4;
  assign wd_fu_1256_p1 = tmp_36_i_fu_1246_p4;
  assign wl_code_table_address0 = tmp_s_fu_566_p1;
  assign wl_code_table_load_c_fu_622_p0 = wl_code_table_q0;
  assign wl_code_table_load_c_fu_622_p1 = wl_code_table_load_c_fu_622_p0;
  assign xd_fu_1819_p2 = (working_key[2224] == 1'b1)? rl_cast_reg_2057 * rh_fu_1801_p2 : rl_cast_reg_2057 - rh_fu_1801_p2;
  assign xs_fu_1824_p2 = (working_key[2225] == 1'b1)? rh_fu_1801_p2 + rl_cast_reg_2057 : rh_fu_1801_p2 - rl_cast_reg_2057;
  assign zl_5_fu_587_p2 = (working_key[2226] == 1'b1)? tmp_i_reg_1928 << zl1_i_reg_378 : tmp_i_reg_1928 + zl1_i_reg_378;
  assign zl_6_fu_1302_p2 = (working_key[2227] == 1'b1)? tmp_i8_33_reg_2096 + zl1_i2_reg_399 : tmp_i8_33_reg_2096 * zl1_i2_reg_399;
  assign zl_fu_499_p2 = (working_key[2228] == 1'b1)? reg_477 - reg_481 : reg_477 * reg_481;
  assign working_key = { locking_key[1873:0] };

endmodule



module backprop_0_obf
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  weights_address0,
  weights_ce0,
  weights_we0,
  weights_d0,
  weights_q0,
  inputs_address0,
  inputs_ce0,
  inputs_q0,
  targets_address0,
  targets_ce0,
  targets_q0,
);

  parameter ap_ST_fsm_state1 = 201'd1;
  parameter ap_ST_fsm_state2 = 201'd2;
  parameter ap_ST_fsm_state3 = 201'd4;
  parameter ap_ST_fsm_state4 = 201'd8;
  parameter ap_ST_fsm_state5 = 201'd16;
  parameter ap_ST_fsm_state6 = 201'd32;
  parameter ap_ST_fsm_state7 = 201'd64;
  parameter ap_ST_fsm_state8 = 201'd128;
  parameter ap_ST_fsm_state9 = 201'd256;
  parameter ap_ST_fsm_state10 = 201'd512;
  parameter ap_ST_fsm_state11 = 201'd1024;
  parameter ap_ST_fsm_state12 = 201'd2048;
  parameter ap_ST_fsm_state13 = 201'd4096;
  parameter ap_ST_fsm_state14 = 201'd8192;
  parameter ap_ST_fsm_state15 = 201'd16384;
  parameter ap_ST_fsm_state16 = 201'd32768;
  parameter ap_ST_fsm_state17 = 201'd65536;
  parameter ap_ST_fsm_state18 = 201'd131072;
  parameter ap_ST_fsm_state19 = 201'd262144;
  parameter ap_ST_fsm_state20 = 201'd524288;
  parameter ap_ST_fsm_state21 = 201'd1048576;
  parameter ap_ST_fsm_state22 = 201'd2097152;
  parameter ap_ST_fsm_state23 = 201'd4194304;
  parameter ap_ST_fsm_state24 = 201'd8388608;
  parameter ap_ST_fsm_state25 = 201'd16777216;
  parameter ap_ST_fsm_state26 = 201'd33554432;
  parameter ap_ST_fsm_state27 = 201'd67108864;
  parameter ap_ST_fsm_state28 = 201'd134217728;
  parameter ap_ST_fsm_state29 = 201'd268435456;
  parameter ap_ST_fsm_state30 = 201'd536870912;
  parameter ap_ST_fsm_state31 = 201'd1073741824;
  parameter ap_ST_fsm_state32 = 201'd2147483648;
  parameter ap_ST_fsm_state33 = 201'd4294967296;
  parameter ap_ST_fsm_state34 = 201'd8589934592;
  parameter ap_ST_fsm_state35 = 201'd17179869184;
  parameter ap_ST_fsm_state36 = 201'd34359738368;
  parameter ap_ST_fsm_state37 = 201'd68719476736;
  parameter ap_ST_fsm_state38 = 201'd137438953472;
  parameter ap_ST_fsm_state39 = 201'd274877906944;
  parameter ap_ST_fsm_state40 = 201'd549755813888;
  parameter ap_ST_fsm_state41 = 201'd1099511627776;
  parameter ap_ST_fsm_state42 = 201'd2199023255552;
  parameter ap_ST_fsm_state43 = 201'd4398046511104;
  parameter ap_ST_fsm_state44 = 201'd8796093022208;
  parameter ap_ST_fsm_state45 = 201'd17592186044416;
  parameter ap_ST_fsm_state46 = 201'd35184372088832;
  parameter ap_ST_fsm_state47 = 201'd70368744177664;
  parameter ap_ST_fsm_state48 = 201'd140737488355328;
  parameter ap_ST_fsm_state49 = 201'd281474976710656;
  parameter ap_ST_fsm_state50 = 201'd562949953421312;
  parameter ap_ST_fsm_state51 = 201'd1125899906842624;
  parameter ap_ST_fsm_state52 = 201'd2251799813685248;
  parameter ap_ST_fsm_state53 = 201'd4503599627370496;
  parameter ap_ST_fsm_state54 = 201'd9007199254740992;
  parameter ap_ST_fsm_state55 = 201'd18014398509481984;
  parameter ap_ST_fsm_state56 = 201'd36028797018963968;
  parameter ap_ST_fsm_state57 = 201'd72057594037927936;
  parameter ap_ST_fsm_state58 = 201'd144115188075855872;
  parameter ap_ST_fsm_state59 = 201'd288230376151711744;
  parameter ap_ST_fsm_state60 = 201'd576460752303423488;
  parameter ap_ST_fsm_state61 = 201'd1152921504606846976;
  parameter ap_ST_fsm_state62 = 201'd2305843009213693952;
  parameter ap_ST_fsm_state63 = 201'd4611686018427387904;
  parameter ap_ST_fsm_state64 = 201'd9223372036854775808;
  parameter ap_ST_fsm_state65 = 201'd18446744073709551616;
  parameter ap_ST_fsm_state66 = 201'd36893488147419103232;
  parameter ap_ST_fsm_state67 = 201'd73786976294838206464;
  parameter ap_ST_fsm_state68 = 201'd147573952589676412928;
  parameter ap_ST_fsm_state69 = 201'd295147905179352825856;
  parameter ap_ST_fsm_state70 = 201'd590295810358705651712;
  parameter ap_ST_fsm_state71 = 201'd1180591620717411303424;
  parameter ap_ST_fsm_state72 = 201'd2361183241434822606848;
  parameter ap_ST_fsm_state73 = 201'd4722366482869645213696;
  parameter ap_ST_fsm_state74 = 201'd9444732965739290427392;
  parameter ap_ST_fsm_state75 = 201'd18889465931478580854784;
  parameter ap_ST_fsm_state76 = 201'd37778931862957161709568;
  parameter ap_ST_fsm_state77 = 201'd75557863725914323419136;
  parameter ap_ST_fsm_state78 = 201'd151115727451828646838272;
  parameter ap_ST_fsm_state79 = 201'd302231454903657293676544;
  parameter ap_ST_fsm_state80 = 201'd604462909807314587353088;
  parameter ap_ST_fsm_state81 = 201'd1208925819614629174706176;
  parameter ap_ST_fsm_state82 = 201'd2417851639229258349412352;
  parameter ap_ST_fsm_state83 = 201'd4835703278458516698824704;
  parameter ap_ST_fsm_state84 = 201'd9671406556917033397649408;
  parameter ap_ST_fsm_state85 = 201'd19342813113834066795298816;
  parameter ap_ST_fsm_state86 = 201'd38685626227668133590597632;
  parameter ap_ST_fsm_state87 = 201'd77371252455336267181195264;
  parameter ap_ST_fsm_state88 = 201'd154742504910672534362390528;
  parameter ap_ST_fsm_state89 = 201'd309485009821345068724781056;
  parameter ap_ST_fsm_state90 = 201'd618970019642690137449562112;
  parameter ap_ST_fsm_state91 = 201'd1237940039285380274899124224;
  parameter ap_ST_fsm_state92 = 201'd2475880078570760549798248448;
  parameter ap_ST_fsm_state93 = 201'd4951760157141521099596496896;
  parameter ap_ST_fsm_state94 = 201'd9903520314283042199192993792;
  parameter ap_ST_fsm_state95 = 201'd19807040628566084398385987584;
  parameter ap_ST_fsm_state96 = 201'd39614081257132168796771975168;
  parameter ap_ST_fsm_state97 = 201'd79228162514264337593543950336;
  parameter ap_ST_fsm_state98 = 201'd158456325028528675187087900672;
  parameter ap_ST_fsm_state99 = 201'd316912650057057350374175801344;
  parameter ap_ST_fsm_state100 = 201'd633825300114114700748351602688;
  parameter ap_ST_fsm_state101 = 201'd1267650600228229401496703205376;
  parameter ap_ST_fsm_state102 = 201'd2535301200456458802993406410752;
  parameter ap_ST_fsm_state103 = 201'd5070602400912917605986812821504;
  parameter ap_ST_fsm_state104 = 201'd10141204801825835211973625643008;
  parameter ap_ST_fsm_state105 = 201'd20282409603651670423947251286016;
  parameter ap_ST_fsm_state106 = 201'd40564819207303340847894502572032;
  parameter ap_ST_fsm_state107 = 201'd81129638414606681695789005144064;
  parameter ap_ST_fsm_state108 = 201'd162259276829213363391578010288128;
  parameter ap_ST_fsm_state109 = 201'd324518553658426726783156020576256;
  parameter ap_ST_fsm_state110 = 201'd649037107316853453566312041152512;
  parameter ap_ST_fsm_state111 = 201'd1298074214633706907132624082305024;
  parameter ap_ST_fsm_state112 = 201'd2596148429267413814265248164610048;
  parameter ap_ST_fsm_state113 = 201'd5192296858534827628530496329220096;
  parameter ap_ST_fsm_state114 = 201'd10384593717069655257060992658440192;
  parameter ap_ST_fsm_state115 = 201'd20769187434139310514121985316880384;
  parameter ap_ST_fsm_state116 = 201'd41538374868278621028243970633760768;
  parameter ap_ST_fsm_state117 = 201'd83076749736557242056487941267521536;
  parameter ap_ST_fsm_state118 = 201'd166153499473114484112975882535043072;
  parameter ap_ST_fsm_state119 = 201'd332306998946228968225951765070086144;
  parameter ap_ST_fsm_state120 = 201'd664613997892457936451903530140172288;
  parameter ap_ST_fsm_state121 = 201'd1329227995784915872903807060280344576;
  parameter ap_ST_fsm_state122 = 201'd2658455991569831745807614120560689152;
  parameter ap_ST_fsm_state123 = 201'd5316911983139663491615228241121378304;
  parameter ap_ST_fsm_state124 = 201'd10633823966279326983230456482242756608;
  parameter ap_ST_fsm_state125 = 201'd21267647932558653966460912964485513216;
  parameter ap_ST_fsm_state126 = 201'd42535295865117307932921825928971026432;
  parameter ap_ST_fsm_state127 = 201'd85070591730234615865843651857942052864;
  parameter ap_ST_fsm_state128 = 201'd170141183460469231731687303715884105728;
  parameter ap_ST_fsm_state129 = 201'd340282366920938463463374607431768211456;
  parameter ap_ST_fsm_state130 = 201'd680564733841876926926749214863536422912;
  parameter ap_ST_fsm_state131 = 201'd1361129467683753853853498429727072845824;
  parameter ap_ST_fsm_state132 = 201'd2722258935367507707706996859454145691648;
  parameter ap_ST_fsm_state133 = 201'd5444517870735015415413993718908291383296;
  parameter ap_ST_fsm_state134 = 201'd10889035741470030830827987437816582766592;
  parameter ap_ST_fsm_state135 = 201'd21778071482940061661655974875633165533184;
  parameter ap_ST_fsm_state136 = 201'd43556142965880123323311949751266331066368;
  parameter ap_ST_fsm_state137 = 201'd87112285931760246646623899502532662132736;
  parameter ap_ST_fsm_state138 = 201'd174224571863520493293247799005065324265472;
  parameter ap_ST_fsm_state139 = 201'd348449143727040986586495598010130648530944;
  parameter ap_ST_fsm_state140 = 201'd696898287454081973172991196020261297061888;
  parameter ap_ST_fsm_state141 = 201'd1393796574908163946345982392040522594123776;
  parameter ap_ST_fsm_state142 = 201'd2787593149816327892691964784081045188247552;
  parameter ap_ST_fsm_state143 = 201'd5575186299632655785383929568162090376495104;
  parameter ap_ST_fsm_state144 = 201'd11150372599265311570767859136324180752990208;
  parameter ap_ST_fsm_state145 = 201'd22300745198530623141535718272648361505980416;
  parameter ap_ST_fsm_state146 = 201'd44601490397061246283071436545296723011960832;
  parameter ap_ST_fsm_state147 = 201'd89202980794122492566142873090593446023921664;
  parameter ap_ST_fsm_state148 = 201'd178405961588244985132285746181186892047843328;
  parameter ap_ST_fsm_state149 = 201'd356811923176489970264571492362373784095686656;
  parameter ap_ST_fsm_state150 = 201'd713623846352979940529142984724747568191373312;
  parameter ap_ST_fsm_state151 = 201'd1427247692705959881058285969449495136382746624;
  parameter ap_ST_fsm_state152 = 201'd2854495385411919762116571938898990272765493248;
  parameter ap_ST_fsm_state153 = 201'd5708990770823839524233143877797980545530986496;
  parameter ap_ST_fsm_state154 = 201'd11417981541647679048466287755595961091061972992;
  parameter ap_ST_fsm_state155 = 201'd22835963083295358096932575511191922182123945984;
  parameter ap_ST_fsm_state156 = 201'd45671926166590716193865151022383844364247891968;
  parameter ap_ST_fsm_state157 = 201'd91343852333181432387730302044767688728495783936;
  parameter ap_ST_fsm_state158 = 201'd182687704666362864775460604089535377456991567872;
  parameter ap_ST_fsm_state159 = 201'd365375409332725729550921208179070754913983135744;
  parameter ap_ST_fsm_state160 = 201'd730750818665451459101842416358141509827966271488;
  parameter ap_ST_fsm_state161 = 201'd1461501637330902918203684832716283019655932542976;
  parameter ap_ST_fsm_state162 = 201'd2923003274661805836407369665432566039311865085952;
  parameter ap_ST_fsm_state163 = 201'd5846006549323611672814739330865132078623730171904;
  parameter ap_ST_fsm_state164 = 201'd11692013098647223345629478661730264157247460343808;
  parameter ap_ST_fsm_state165 = 201'd23384026197294446691258957323460528314494920687616;
  parameter ap_ST_fsm_state166 = 201'd46768052394588893382517914646921056628989841375232;
  parameter ap_ST_fsm_state167 = 201'd93536104789177786765035829293842113257979682750464;
  parameter ap_ST_fsm_state168 = 201'd187072209578355573530071658587684226515959365500928;
  parameter ap_ST_fsm_state169 = 201'd374144419156711147060143317175368453031918731001856;
  parameter ap_ST_fsm_state170 = 201'd748288838313422294120286634350736906063837462003712;
  parameter ap_ST_fsm_state171 = 201'd1496577676626844588240573268701473812127674924007424;
  parameter ap_ST_fsm_state172 = 201'd2993155353253689176481146537402947624255349848014848;
  parameter ap_ST_fsm_state173 = 201'd5986310706507378352962293074805895248510699696029696;
  parameter ap_ST_fsm_state174 = 201'd11972621413014756705924586149611790497021399392059392;
  parameter ap_ST_fsm_state175 = 201'd23945242826029513411849172299223580994042798784118784;
  parameter ap_ST_fsm_state176 = 201'd47890485652059026823698344598447161988085597568237568;
  parameter ap_ST_fsm_state177 = 201'd95780971304118053647396689196894323976171195136475136;
  parameter ap_ST_fsm_state178 = 201'd191561942608236107294793378393788647952342390272950272;
  parameter ap_ST_fsm_state179 = 201'd383123885216472214589586756787577295904684780545900544;
  parameter ap_ST_fsm_state180 = 201'd766247770432944429179173513575154591809369561091801088;
  parameter ap_ST_fsm_state181 = 201'd1532495540865888858358347027150309183618739122183602176;
  parameter ap_ST_fsm_state182 = 201'd3064991081731777716716694054300618367237478244367204352;
  parameter ap_ST_fsm_state183 = 201'd6129982163463555433433388108601236734474956488734408704;
  parameter ap_ST_fsm_state184 = 201'd12259964326927110866866776217202473468949912977468817408;
  parameter ap_ST_fsm_state185 = 201'd24519928653854221733733552434404946937899825954937634816;
  parameter ap_ST_fsm_state186 = 201'd49039857307708443467467104868809893875799651909875269632;
  parameter ap_ST_fsm_state187 = 201'd98079714615416886934934209737619787751599303819750539264;
  parameter ap_ST_fsm_state188 = 201'd196159429230833773869868419475239575503198607639501078528;
  parameter ap_ST_fsm_state189 = 201'd392318858461667547739736838950479151006397215279002157056;
  parameter ap_ST_fsm_state190 = 201'd784637716923335095479473677900958302012794430558004314112;
  parameter ap_ST_fsm_state191 = 201'd1569275433846670190958947355801916604025588861116008628224;
  parameter ap_ST_fsm_state192 = 201'd3138550867693340381917894711603833208051177722232017256448;
  parameter ap_ST_fsm_state193 = 201'd6277101735386680763835789423207666416102355444464034512896;
  parameter ap_ST_fsm_state194 = 201'd12554203470773361527671578846415332832204710888928069025792;
  parameter ap_ST_fsm_state195 = 201'd25108406941546723055343157692830665664409421777856138051584;
  parameter ap_ST_fsm_state196 = 201'd50216813883093446110686315385661331328818843555712276103168;
  parameter ap_ST_fsm_state197 = 201'd100433627766186892221372630771322662657637687111424552206336;
  parameter ap_ST_fsm_state198 = 201'd200867255532373784442745261542645325315275374222849104412672;
  parameter ap_ST_fsm_state199 = 201'd401734511064747568885490523085290650630550748445698208825344;
  parameter ap_ST_fsm_state200 = 201'd803469022129495137770981046170581301261101496891396417650688;
  parameter ap_ST_fsm_state201 = 201'd1606938044258990275541962092341162602522202993782792835301376;
  input ap_clk;
  input ap_rst;
  input ap_start;
  input [39:0] working_key;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [7:0] weights_address0;
  output weights_ce0;
  output weights_we0;
  output [63:0] weights_d0;
  input [63:0] weights_q0;
  output [8:0] inputs_address0;
  output inputs_ce0;
  input [63:0] inputs_q0;
  output [9:0] targets_address0;
  output targets_ce0;
  input [63:0] targets_q0;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [7:0] weights_address0;
  reg weights_ce0;
  reg weights_we0;
  reg inputs_ce0;
  reg targets_ce0;
  reg [200:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  wire [63:0] activations_q0;
  reg [63:0] reg_583;
  wire ap_CS_fsm_state14;
  wire ap_CS_fsm_state69;
  wire ap_CS_fsm_state178;
  reg [63:0] reg_590;
  wire ap_CS_fsm_state118;
  wire ap_CS_fsm_state190;
  wire [63:0] grp_fu_566_p2;
  reg [63:0] reg_596;
  wire ap_CS_fsm_state19;
  wire ap_CS_fsm_state114;
  wire ap_CS_fsm_state123;
  wire ap_CS_fsm_state174;
  wire ap_CS_fsm_state185;
  wire ap_CS_fsm_state195;
  wire [63:0] grp_fu_578_p2;
  reg [63:0] reg_604;
  wire ap_CS_fsm_state37;
  wire ap_CS_fsm_state82;
  wire ap_CS_fsm_state142;
  wire [63:0] grp_fu_559_p2;
  reg [63:0] reg_609;
  wire ap_CS_fsm_state42;
  wire ap_CS_fsm_state74;
  wire ap_CS_fsm_state147;
  wire ap_CS_fsm_state200;
  wire [63:0] grp_fu_573_p2;
  reg [63:0] reg_617;
  wire ap_CS_fsm_state64;
  wire ap_CS_fsm_state109;
  wire ap_CS_fsm_state169;
  wire [63:0] deltas_q0;
  reg [63:0] reg_623;
  wire ap_CS_fsm_state180;
  wire [1:0] ee_fu_634_p2;
  reg [1:0] ee_reg_1581;
  wire ap_CS_fsm_state2;
  wire [5:0] add_ln160_fu_664_p2;
  reg [5:0] add_ln160_reg_1586;
  wire [0:0] icmp_ln156_fu_628_p2;
  wire [3:0] rows_fu_676_p2;
  reg [3:0] rows_reg_1594;
  wire ap_CS_fsm_state3;
  wire [9:0] add_ln160_2_fu_720_p2;
  reg [9:0] add_ln160_2_reg_1599;
  wire [0:0] icmp_ln157_fu_670_p2;
  wire [3:0] cols_fu_732_p2;
  wire ap_CS_fsm_state4;
  wire [6:0] ee_2_fu_758_p2;
  reg [6:0] ee_2_reg_1615;
  wire ap_CS_fsm_state5;
  wire [6:0] jj_1_fu_770_p2;
  reg [6:0] jj_1_reg_1623;
  wire ap_CS_fsm_state6;
  wire [1:0] cols_2_fu_782_p2;
  reg [1:0] cols_2_reg_1631;
  wire ap_CS_fsm_state7;
  wire [5:0] add_ln170_fu_812_p2;
  reg [5:0] add_ln170_reg_1636;
  wire [0:0] icmp_ln168_fu_776_p2;
  wire [9:0] zext_ln52_fu_826_p1;
  reg [9:0] zext_ln52_reg_1641;
  wire [10:0] add_ln52_fu_854_p2;
  reg [10:0] add_ln52_reg_1646;
  wire [3:0] rows_2_fu_866_p2;
  wire ap_CS_fsm_state8;
  wire [2:0] i_fu_892_p2;
  reg [2:0] i_reg_1662;
  wire ap_CS_fsm_state9;
  wire [0:0] icmp_ln34_fu_886_p2;
  wire [1:0] i_1_fu_923_p2;
  reg [1:0] i_1_reg_1675;
  wire ap_CS_fsm_state11;
  wire [5:0] add_ln21_fu_953_p2;
  reg [5:0] add_ln21_reg_1680;
  wire [0:0] icmp_ln39_fu_917_p2;
  wire [3:0] select_ln40_fu_963_p3;
  reg [3:0] select_ln40_reg_1685;
  wire [5:0] add_ln23_fu_995_p2;
  reg [5:0] add_ln23_reg_1690;
  wire [3:0] ii_fu_1007_p2;
  reg [3:0] ii_reg_1698;
  wire ap_CS_fsm_state12;
  wire [8:0] zext_ln23_2_fu_1013_p1;
  reg [8:0] zext_ln23_2_reg_1703;
  wire [0:0] icmp_ln18_fu_1001_p2;
  reg [4:0] activations_addr_5_reg_1708;
  wire [3:0] jj_fu_1036_p2;
  reg [3:0] jj_reg_1716;
  wire ap_CS_fsm_state13;
  wire [0:0] icmp_ln20_fu_1031_p2;
  wire [63:0] xor_ln7_1_fu_1096_p2;
  reg [63:0] xor_ln7_1_reg_1731;
  wire ap_CS_fsm_state24;
  wire [63:0] bitcast_ln7_3_fu_1102_p1;
  wire ap_CS_fsm_state25;
  wire [1:0] i_3_fu_1112_p2;
  reg [1:0] i_3_reg_1749;
  wire ap_CS_fsm_state66;
  wire [5:0] add_ln112_fu_1142_p2;
  reg [5:0] add_ln112_reg_1754;
  wire [0:0] icmp_ln110_fu_1106_p2;
  wire [3:0] j_fu_1154_p2;
  wire ap_CS_fsm_state67;
  wire [3:0] i_2_fu_1180_p2;
  reg [3:0] i_2_reg_1770;
  wire ap_CS_fsm_state68;
  wire [4:0] zext_ln52_3_fu_1186_p1;
  reg [4:0] zext_ln52_3_reg_1775;
  wire [0:0] icmp_ln51_fu_1174_p2;
  reg [63:0] targets_load_reg_1790;
  wire [63:0] xor_ln7_fu_1219_p2;
  reg [63:0] xor_ln7_reg_1795;
  wire [63:0] bitcast_ln7_1_fu_1225_p1;
  wire ap_CS_fsm_state70;
  reg [63:0] temp_reg_1805;
  wire ap_CS_fsm_state87;
  wire [3:0] add_ln70_fu_1245_p2;
  reg [3:0] add_ln70_reg_1813;
  wire ap_CS_fsm_state116;
  wire [8:0] add_ln73_1_fu_1295_p2;
  reg [8:0] add_ln73_1_reg_1818;
  wire [0:0] icmp_ln70_fu_1239_p2;
  reg [4:0] deltas_addr_2_reg_1823;
  reg [4:0] activations_addr_6_reg_1828;
  wire [3:0] add_ln72_fu_1307_p2;
  reg [3:0] add_ln72_reg_1836;
  wire ap_CS_fsm_state117;
  wire [0:0] icmp_ln72_fu_1301_p2;
  wire ap_CS_fsm_state128;
  wire [63:0] xor_ln7_2_fu_1346_p2;
  reg [63:0] xor_ln7_2_reg_1856;
  wire ap_CS_fsm_state129;
  wire [63:0] bitcast_ln7_5_fu_1352_p1;
  wire ap_CS_fsm_state130;
  wire [1:0] j_2_fu_1362_p2;
  reg [1:0] j_2_reg_1869;
  wire ap_CS_fsm_state176;
  wire [0:0] icmp_ln123_fu_1356_p2;
  wire [5:0] add_ln90_fu_1392_p2;
  reg [5:0] add_ln90_reg_1874;
  wire [5:0] add_ln90_1_fu_1422_p2;
  reg [5:0] add_ln90_1_reg_1880;
  wire [3:0] select_ln87_fu_1434_p3;
  reg [3:0] select_ln87_reg_1885;
  wire [3:0] ii_1_fu_1447_p2;
  reg [3:0] ii_1_reg_1893;
  wire ap_CS_fsm_state177;
  wire [5:0] add_ln90_2_fu_1457_p2;
  reg [5:0] add_ln90_2_reg_1898;
  wire [0:0] icmp_ln87_fu_1442_p2;
  wire [5:0] add_ln90_4_fu_1467_p2;
  reg [5:0] add_ln90_4_reg_1904;
  wire [8:0] add_ln90_3_fu_1490_p2;
  reg [8:0] add_ln90_3_reg_1915;
  wire [9:0] add_ln90_5_fu_1518_p2;
  reg [9:0] add_ln90_5_reg_1920;
  wire [3:0] jj_2_fu_1530_p2;
  reg [3:0] jj_2_reg_1928;
  wire ap_CS_fsm_state179;
  reg [7:0] weights_addr_2_reg_1933;
  wire [0:0] icmp_ln88_fu_1524_p2;
  reg [8:0] changeMat_addr_1_reg_1943;
  wire [63:0] changeMat_q0;
  reg [63:0] changeMat_load_reg_1948;
  wire ap_CS_fsm_state187;
  reg [4:0] deltas_address0;
  reg deltas_ce0;
  reg deltas_we0;
  reg [63:0] deltas_d0;
  reg [8:0] changeMat_address0;
  reg changeMat_ce0;
  reg changeMat_we0;
  reg [63:0] changeMat_d0;
  reg [4:0] activations_address0;
  reg activations_ce0;
  reg activations_we0;
  reg [63:0] activations_d0;
  reg [1:0] ee_0_reg_324;
  reg [3:0] rows_0_reg_335;
  wire [0:0] icmp_ln159_fu_726_p2;
  reg [3:0] cols_0_reg_346;
  reg [6:0] ee_1_reg_357;
  wire [0:0] icmp_ln167_fu_764_p2;
  reg [6:0] jj_0_reg_368;
  wire [0:0] icmp_ln165_fu_752_p2;
  reg [1:0] cols_1_reg_380;
  wire [0:0] icmp_ln169_fu_860_p2;
  reg [3:0] rows_1_reg_391;
  reg [2:0] i_0_i_reg_402;
  wire ap_CS_fsm_state10;
  reg [1:0] i_1_i_reg_414;
  reg [3:0] ii_0_i_i_reg_425;
  wire ap_CS_fsm_state65;
  reg [3:0] jj_0_i_i_reg_436;
  reg [63:0] x_assign_1_reg_447;
  reg [1:0] i_0_i13_reg_459;
  wire [0:0] icmp_ln111_fu_1148_p2;
  reg [3:0] j_0_i_reg_470;
  reg [3:0] i_0_i_i_reg_481;
  wire ap_CS_fsm_state115;
  reg [3:0] jj_0_i_i21_0_reg_492;
  wire ap_CS_fsm_state175;
  reg [3:0] kk_0_i_i_0_reg_503;
  reg [63:0] error_0_i_i_0_reg_514;
  reg [1:0] level_assign_reg_526;
  reg [3:0] ii_0_i_i25_reg_537;
  reg [3:0] jj_0_i10_i_reg_548;
  wire ap_CS_fsm_state201;
  wire [63:0] zext_ln160_3_fu_691_p1;
  wire [63:0] zext_ln160_7_fu_747_p1;
  wire [63:0] zext_ln170_3_fu_881_p1;
  wire [63:0] zext_ln35_2_fu_907_p1;
  wire [63:0] zext_ln35_fu_912_p1;
  wire [63:0] zext_ln23_4_fu_1026_p1;
  wire [63:0] zext_ln21_5_fu_1087_p1;
  wire [63:0] zext_ln21_3_fu_1051_p1;
  wire [63:0] zext_ln112_3_fu_1169_p1;
  wire [63:0] zext_ln52_5_fu_1199_p1;
  wire [63:0] zext_ln52_6_fu_1210_p1;
  wire [63:0] zext_ln53_fu_1234_p1;
  wire [63:0] zext_ln73_fu_1251_p1;
  wire [63:0] zext_ln73_2_fu_1266_p1;
  wire [63:0] zext_ln73_7_fu_1326_p1;
  wire [63:0] zext_ln73_8_fu_1337_p1;
  wire [63:0] zext_ln90_5_fu_1462_p1;
  wire [63:0] zext_ln90_12_fu_1553_p1;
  wire [63:0] zext_ln89_fu_1563_p1;
  wire [63:0] zext_ln90_13_fu_1573_p1;
  wire ap_CS_fsm_state186;
  wire ap_CS_fsm_state189;
  reg [63:0] grp_fu_559_p0;
  reg [63:0] grp_fu_559_p1;
  wire ap_CS_fsm_state20;
  wire ap_CS_fsm_state38;
  wire ap_CS_fsm_state83;
  wire ap_CS_fsm_state124;
  wire ap_CS_fsm_state143;
  wire ap_CS_fsm_state191;
  wire ap_CS_fsm_state196;
  reg [63:0] grp_fu_566_p0;
  reg [63:0] grp_fu_566_p1;
  wire ap_CS_fsm_state15;
  wire ap_CS_fsm_state110;
  wire ap_CS_fsm_state119;
  wire ap_CS_fsm_state170;
  wire ap_CS_fsm_state181;
  reg [63:0] grp_fu_573_p1;
  wire ap_CS_fsm_state43;
  wire ap_CS_fsm_state88;
  wire ap_CS_fsm_state148;
  reg [63:0] grp_fu_578_p1;
  wire [4:0] tmp_fu_640_p3;
  wire [2:0] tmp_19_fu_652_p3;
  wire [5:0] zext_ln160_1_fu_660_p1;
  wire [5:0] zext_ln160_fu_648_p1;
  wire [5:0] zext_ln160_2_fu_682_p1;
  wire [5:0] add_ln160_1_fu_686_p2;
  wire [8:0] tmp_20_fu_696_p3;
  wire [6:0] tmp_21_fu_708_p3;
  wire [9:0] zext_ln160_4_fu_704_p1;
  wire [9:0] zext_ln160_5_fu_716_p1;
  wire [9:0] zext_ln160_6_fu_738_p1;
  wire [9:0] add_ln160_3_fu_742_p2;
  wire [4:0] tmp_25_fu_788_p3;
  wire [2:0] tmp_26_fu_800_p3;
  wire [5:0] zext_ln170_1_fu_808_p1;
  wire [5:0] zext_ln170_fu_796_p1;
  wire [8:0] tmp_22_fu_818_p3;
  wire [9:0] tmp_23_fu_830_p3;
  wire [7:0] tmp_24_fu_842_p3;
  wire [10:0] zext_ln52_2_fu_850_p1;
  wire [10:0] zext_ln52_1_fu_838_p1;
  wire [5:0] zext_ln170_2_fu_872_p1;
  wire [5:0] add_ln170_1_fu_876_p2;
  wire [9:0] zext_ln35_1_fu_898_p1;
  wire [9:0] add_ln35_fu_902_p2;
  wire [4:0] tmp_27_fu_929_p3;
  wire [2:0] tmp_28_fu_941_p3;
  wire [5:0] zext_ln21_fu_937_p1;
  wire [5:0] zext_ln21_1_fu_949_p1;
  wire [0:0] trunc_ln40_fu_959_p1;
  wire [4:0] tmp_29_fu_971_p3;
  wire [2:0] tmp_30_fu_983_p3;
  wire [5:0] zext_ln23_fu_979_p1;
  wire [5:0] zext_ln23_1_fu_991_p1;
  wire [5:0] zext_ln23_3_fu_1017_p1;
  wire [5:0] add_ln23_1_fu_1021_p2;
  wire [5:0] zext_ln21_2_fu_1042_p1;
  wire [5:0] add_ln21_1_fu_1046_p2;
  wire [6:0] tmp_33_fu_1064_p3;
  wire [8:0] p_shl_cast_fu_1056_p3;
  wire [8:0] zext_ln21_4_fu_1072_p1;
  wire [8:0] add_ln21_2_fu_1076_p2;
  wire [8:0] add_ln21_3_fu_1082_p2;
  wire [63:0] bitcast_ln7_2_fu_1092_p1;
  wire [4:0] tmp_31_fu_1118_p3;
  wire [2:0] tmp_32_fu_1130_p3;
  wire [5:0] zext_ln112_1_fu_1138_p1;
  wire [5:0] zext_ln112_fu_1126_p1;
  wire [5:0] zext_ln112_2_fu_1160_p1;
  wire [5:0] add_ln112_1_fu_1164_p2;
  wire [10:0] zext_ln52_4_fu_1190_p1;
  wire [10:0] add_ln52_1_fu_1194_p2;
  wire [4:0] add_ln52_2_fu_1204_p2;
  wire [63:0] bitcast_ln7_fu_1215_p1;
  wire [4:0] add_ln53_fu_1229_p2;
  wire [4:0] zext_ln73_1_fu_1256_p1;
  wire [4:0] add_ln73_fu_1260_p2;
  wire [7:0] tmp_34_fu_1271_p3;
  wire [5:0] tmp_35_fu_1283_p3;
  wire [8:0] zext_ln73_3_fu_1279_p1;
  wire [8:0] zext_ln73_4_fu_1291_p1;
  wire [8:0] zext_ln73_6_fu_1317_p1;
  wire [8:0] add_ln73_2_fu_1321_p2;
  wire [4:0] zext_ln73_5_fu_1313_p1;
  wire [4:0] add_ln73_3_fu_1331_p2;
  wire [63:0] bitcast_ln7_4_fu_1342_p1;
  wire [4:0] tmp_36_fu_1368_p3;
  wire [2:0] tmp_37_fu_1380_p3;
  wire [5:0] zext_ln90_1_fu_1388_p1;
  wire [5:0] zext_ln90_fu_1376_p1;
  wire [4:0] tmp_38_fu_1398_p3;
  wire [2:0] tmp_39_fu_1410_p3;
  wire [5:0] zext_ln90_3_fu_1418_p1;
  wire [5:0] zext_ln90_2_fu_1406_p1;
  wire [0:0] icmp_ln87_1_fu_1428_p2;
  wire [5:0] zext_ln90_4_fu_1453_p1;
  wire [6:0] tmp_40_fu_1479_p3;
  wire [8:0] p_shl6_cast_fu_1472_p3;
  wire [8:0] zext_ln90_6_fu_1486_p1;
  wire [8:0] tmp_41_fu_1496_p3;
  wire [6:0] tmp_42_fu_1507_p3;
  wire [9:0] zext_ln90_7_fu_1503_p1;
  wire [9:0] zext_ln90_8_fu_1514_p1;
  wire [8:0] zext_ln90_11_fu_1544_p1;
  wire [8:0] add_ln90_6_fu_1548_p2;
  wire [5:0] zext_ln90_10_fu_1540_p1;
  wire [5:0] add_ln89_fu_1558_p2;
  wire [9:0] zext_ln90_9_fu_1536_p1;
  wire [9:0] add_ln90_7_fu_1568_p2;
  reg [1:0] grp_fu_559_opcode;
  reg [200:0] ap_NS_fsm;

  initial begin
    #0 ap_CS_fsm = 201'd1;
  end


  backprop_deltas
  #(
    .DataWidth(64),
    .AddressRange(30),
    .AddressWidth(5)
  )
  deltas_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(deltas_address0),
    .ce0(deltas_ce0),
    .we0(deltas_we0),
    .d0(deltas_d0),
    .q0(deltas_q0)
  );


  backprop_changeMat
  #(
    .DataWidth(64),
    .AddressRange(300),
    .AddressWidth(9)
  )
  changeMat_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(changeMat_address0),
    .ce0(changeMat_ce0),
    .we0(changeMat_we0),
    .d0(changeMat_d0),
    .q0(changeMat_q0)
  );


  backprop_deltas
  #(
    .DataWidth(64),
    .AddressRange(30),
    .AddressWidth(5)
  )
  activations_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(activations_address0),
    .ce0(activations_ce0),
    .we0(activations_we0),
    .d0(activations_d0),
    .q0(activations_q0)
  );


  backprop_dadddsubcud
  #(
    .ID(1),
    .NUM_STAGE(5),
    .din0_WIDTH(64),
    .din1_WIDTH(64),
    .dout_WIDTH(64)
  )
  backprop_dadddsubcud_U1
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_559_p0),
    .din1(grp_fu_559_p1),
    .opcode(grp_fu_559_opcode),
    .ce(1'b1),
    .dout(grp_fu_559_p2)
  );


  backprop_dmul_64ndEe
  #(
    .ID(1),
    .NUM_STAGE(5),
    .din0_WIDTH(64),
    .din1_WIDTH(64),
    .dout_WIDTH(64)
  )
  backprop_dmul_64ndEe_U2
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_566_p0),
    .din1(grp_fu_566_p1),
    .ce(1'b1),
    .dout(grp_fu_566_p2)
  );


  backprop_ddiv_64neOg
  #(
    .ID(1),
    .NUM_STAGE(22),
    .din0_WIDTH(64),
    .din1_WIDTH(64),
    .dout_WIDTH(64)
  )
  backprop_ddiv_64neOg_U3
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(64'd4607182418800017408),
    .din1(grp_fu_573_p1),
    .ce(1'b1),
    .dout(grp_fu_573_p2)
  );


  backprop_dexp_64nfYi
  #(
    .ID(1),
    .NUM_STAGE(13),
    .din0_WIDTH(64),
    .din1_WIDTH(64),
    .dout_WIDTH(64)
  )
  backprop_dexp_64nfYi_U4
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(64'd0),
    .din1(grp_fu_578_p1),
    .ce(1'b1),
    .dout(grp_fu_578_p2)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if((icmp_ln159_fu_726_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state4)) begin
      cols_0_reg_346 <= cols_fu_732_p2;
    end else if((icmp_ln157_fu_670_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3)) begin
      cols_0_reg_346 <= 4'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln169_fu_860_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state8)) begin
      cols_1_reg_380 <= cols_2_reg_1631;
    end else if((icmp_ln167_fu_764_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state6)) begin
      cols_1_reg_380 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln157_fu_670_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state3)) begin
      ee_0_reg_324 <= ee_reg_1581;
    end else if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      ee_0_reg_324 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln156_fu_628_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
      ee_1_reg_357 <= 7'd0;
    end else if((icmp_ln167_fu_764_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state6)) begin
      ee_1_reg_357 <= ee_2_reg_1615;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state128) begin
      error_0_i_i_0_reg_514 <= grp_fu_559_p2;
    end else if((icmp_ln70_fu_1239_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state116)) begin
      error_0_i_i_0_reg_514 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln39_fu_917_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state11)) begin
      i_0_i13_reg_459 <= 2'd0;
    end else if((icmp_ln111_fu_1148_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state67)) begin
      i_0_i13_reg_459 <= i_3_reg_1749;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln110_fu_1106_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state66)) begin
      i_0_i_i_reg_481 <= 4'd0;
    end else if(1'b1 == ap_CS_fsm_state115) begin
      i_0_i_i_reg_481 <= i_2_reg_1770;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state10) begin
      i_0_i_reg_402 <= i_reg_1662;
    end else if((icmp_ln168_fu_776_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state7)) begin
      i_0_i_reg_402 <= 3'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln34_fu_886_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state9)) begin
      i_1_i_reg_414 <= 2'd0;
    end else if((icmp_ln18_fu_1001_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state12)) begin
      i_1_i_reg_414 <= i_1_reg_1675;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln88_fu_1524_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state179)) begin
      ii_0_i_i25_reg_537 <= ii_1_reg_1893;
    end else if((icmp_ln123_fu_1356_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state176)) begin
      ii_0_i_i25_reg_537 <= 4'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state65) begin
      ii_0_i_i_reg_425 <= ii_reg_1698;
    end else if((icmp_ln39_fu_917_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state11)) begin
      ii_0_i_i_reg_425 <= 4'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln111_fu_1148_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state67)) begin
      j_0_i_reg_470 <= j_fu_1154_p2;
    end else if((icmp_ln110_fu_1106_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state66)) begin
      j_0_i_reg_470 <= 4'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state201) begin
      jj_0_i10_i_reg_548 <= jj_2_reg_1928;
    end else if(1'b1 == ap_CS_fsm_state178) begin
      jj_0_i10_i_reg_548 <= 4'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state175) begin
      jj_0_i_i21_0_reg_492 <= add_ln70_reg_1813;
    end else if((icmp_ln51_fu_1174_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state68)) begin
      jj_0_i_i21_0_reg_492 <= 4'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state24) begin
      jj_0_i_i_reg_436 <= jj_reg_1716;
    end else if((icmp_ln18_fu_1001_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state12)) begin
      jj_0_i_i_reg_436 <= 4'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln123_fu_1356_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state176)) begin
      jj_0_reg_368 <= jj_1_reg_1623;
    end else if((icmp_ln165_fu_752_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state5)) begin
      jj_0_reg_368 <= 7'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state128) begin
      kk_0_i_i_0_reg_503 <= add_ln72_reg_1836;
    end else if((icmp_ln70_fu_1239_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state116)) begin
      kk_0_i_i_0_reg_503 <= 4'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln70_fu_1239_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state116)) begin
      level_assign_reg_526 <= 2'd2;
    end else if((icmp_ln87_fu_1442_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state177)) begin
      level_assign_reg_526 <= j_2_reg_1869;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln159_fu_726_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state4)) begin
      rows_0_reg_335 <= rows_reg_1594;
    end else if((icmp_ln156_fu_628_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      rows_0_reg_335 <= 4'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln169_fu_860_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state8)) begin
      rows_1_reg_391 <= rows_2_fu_866_p2;
    end else if((icmp_ln168_fu_776_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      rows_1_reg_391 <= 4'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state24) begin
      x_assign_1_reg_447 <= grp_fu_559_p2;
    end else if((icmp_ln18_fu_1001_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state12)) begin
      x_assign_1_reg_447 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln18_fu_1001_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state12)) begin
      activations_addr_5_reg_1708 <= zext_ln23_4_fu_1026_p1;
      zext_ln23_2_reg_1703[3:0] <= zext_ln23_2_fu_1013_p1[3:0];
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln70_fu_1239_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state116)) begin
      activations_addr_6_reg_1828 <= zext_ln73_2_fu_1266_p1;
      add_ln73_1_reg_1818[8:1] <= add_ln73_1_fu_1295_p2[8:1];
      deltas_addr_2_reg_1823[3:0] <= zext_ln73_fu_1251_p1[3:0];
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln110_fu_1106_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state66)) begin
      add_ln112_reg_1754[5:1] <= add_ln112_fu_1142_p2[5:1];
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln157_fu_670_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3)) begin
      add_ln160_2_reg_1599[9:1] <= add_ln160_2_fu_720_p2[9:1];
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln156_fu_628_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      add_ln160_reg_1586[5:1] <= add_ln160_fu_664_p2[5:1];
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln168_fu_776_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      add_ln170_reg_1636[5:1] <= add_ln170_fu_812_p2[5:1];
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln39_fu_917_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state11)) begin
      add_ln21_reg_1680[5:1] <= add_ln21_fu_953_p2[5:1];
      add_ln23_reg_1690[5:1] <= add_ln23_fu_995_p2[5:1];
      select_ln40_reg_1685[3:1] <= select_ln40_fu_963_p3[3:1];
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln168_fu_776_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state7)) begin
      add_ln52_reg_1646[10:1] <= add_ln52_fu_854_p2[10:1];
      zext_ln52_reg_1641[8:2] <= zext_ln52_fu_826_p1[8:2];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state116) begin
      add_ln70_reg_1813 <= add_ln70_fu_1245_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state117) begin
      add_ln72_reg_1836 <= add_ln72_fu_1307_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln123_fu_1356_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state176)) begin
      add_ln90_1_reg_1880[5:1] <= add_ln90_1_fu_1422_p2[5:1];
      add_ln90_reg_1874[5:1] <= add_ln90_fu_1392_p2[5:1];
      j_2_reg_1869 <= j_2_fu_1362_p2;
      select_ln87_reg_1885[3:1] <= select_ln87_fu_1434_p3[3:1];
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln87_fu_1442_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state177)) begin
      add_ln90_2_reg_1898 <= add_ln90_2_fu_1457_p2;
      add_ln90_4_reg_1904 <= add_ln90_4_fu_1467_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state178) begin
      add_ln90_3_reg_1915[8:1] <= add_ln90_3_fu_1490_p2[8:1];
      add_ln90_5_reg_1920[9:1] <= add_ln90_5_fu_1518_p2[9:1];
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln88_fu_1524_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state179)) begin
      changeMat_addr_1_reg_1943 <= zext_ln90_13_fu_1573_p1;
      weights_addr_2_reg_1933 <= zext_ln90_12_fu_1553_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state187) begin
      changeMat_load_reg_1948 <= changeMat_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      cols_2_reg_1631 <= cols_2_fu_782_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      ee_2_reg_1615 <= ee_2_fu_758_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      ee_reg_1581 <= ee_fu_634_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      i_1_reg_1675 <= i_1_fu_923_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state68) begin
      i_2_reg_1770 <= i_2_fu_1180_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state66) begin
      i_3_reg_1749 <= i_3_fu_1112_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      i_reg_1662 <= i_fu_892_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state177) begin
      ii_1_reg_1893 <= ii_1_fu_1447_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      ii_reg_1698 <= ii_fu_1007_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state6) begin
      jj_1_reg_1623 <= jj_1_fu_770_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state179) begin
      jj_2_reg_1928 <= jj_2_fu_1530_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      jj_reg_1716 <= jj_fu_1036_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state178) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state14)) begin
      reg_583 <= activations_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state190) | (1'b1 == ap_CS_fsm_state118) | (1'b1 == ap_CS_fsm_state14)) begin
      reg_590 <= weights_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state195) | (1'b1 == ap_CS_fsm_state185) | (1'b1 == ap_CS_fsm_state174) | (1'b1 == ap_CS_fsm_state123) | (1'b1 == ap_CS_fsm_state114) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state190)) begin
      reg_596 <= grp_fu_566_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state142) | (1'b1 == ap_CS_fsm_state82) | (1'b1 == ap_CS_fsm_state37)) begin
      reg_604 <= grp_fu_578_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state200) | (1'b1 == ap_CS_fsm_state147) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state42) | (1'b1 == ap_CS_fsm_state195)) begin
      reg_609 <= grp_fu_559_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state169) | (1'b1 == ap_CS_fsm_state109) | (1'b1 == ap_CS_fsm_state64)) begin
      reg_617 <= grp_fu_573_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state180) | (1'b1 == ap_CS_fsm_state118)) begin
      reg_623 <= deltas_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      rows_reg_1594 <= rows_fu_676_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state69) begin
      targets_load_reg_1790 <= targets_q0;
      xor_ln7_reg_1795 <= xor_ln7_fu_1219_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state87) begin
      temp_reg_1805 <= grp_fu_559_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln20_fu_1031_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state13)) begin
      xor_ln7_1_reg_1731 <= xor_ln7_1_fu_1096_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state129) begin
      xor_ln7_2_reg_1856 <= xor_ln7_2_fu_1346_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln51_fu_1174_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state68)) begin
      zext_ln52_3_reg_1775[3:0] <= zext_ln52_3_fu_1186_p1[3:0];
    end 
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state177) begin
      activations_address0 = zext_ln90_5_fu_1462_p1;
    end else if(1'b1 == ap_CS_fsm_state117) begin
      activations_address0 = activations_addr_6_reg_1828;
    end else if(1'b1 == ap_CS_fsm_state68) begin
      activations_address0 = zext_ln52_6_fu_1210_p1;
    end else if(1'b1 == ap_CS_fsm_state65) begin
      activations_address0 = activations_addr_5_reg_1708;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      activations_address0 = zext_ln21_3_fu_1051_p1;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      activations_address0 = zext_ln35_fu_912_p1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      activations_address0 = zext_ln170_3_fu_881_p1;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      activations_address0 = zext_ln160_3_fu_691_p1;
    end else begin
      activations_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state65) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state177) | (1'b1 == ap_CS_fsm_state117) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state3)) begin
      activations_ce0 = 1'b1;
    end else begin
      activations_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state65) begin
      activations_d0 = reg_617;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      activations_d0 = inputs_q0;
    end else if((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state3)) begin
      activations_d0 = 64'd4607182418800017408;
    end else begin
      activations_d0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state65) | (1'b1 == ap_CS_fsm_state10) | (icmp_ln169_fu_860_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state8) | (icmp_ln157_fu_670_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3)) begin
      activations_we0 = 1'b1;
    end else begin
      activations_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((icmp_ln165_fu_752_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state5)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if((icmp_ln165_fu_752_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state5)) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state186) begin
      changeMat_address0 = changeMat_addr_1_reg_1943;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      changeMat_address0 = zext_ln160_7_fu_747_p1;
    end else begin
      changeMat_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state186) | (1'b1 == ap_CS_fsm_state4)) begin
      changeMat_ce0 = 1'b1;
    end else begin
      changeMat_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state186) begin
      changeMat_d0 = reg_596;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      changeMat_d0 = 64'd0;
    end else begin
      changeMat_d0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state186) | (icmp_ln159_fu_726_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state4)) begin
      changeMat_we0 = 1'b1;
    end else begin
      changeMat_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state179) begin
      deltas_address0 = zext_ln89_fu_1563_p1;
    end else if(1'b1 == ap_CS_fsm_state175) begin
      deltas_address0 = deltas_addr_2_reg_1823;
    end else if(1'b1 == ap_CS_fsm_state117) begin
      deltas_address0 = zext_ln73_8_fu_1337_p1;
    end else if(1'b1 == ap_CS_fsm_state115) begin
      deltas_address0 = zext_ln53_fu_1234_p1;
    end else if(1'b1 == ap_CS_fsm_state67) begin
      deltas_address0 = zext_ln112_3_fu_1169_p1;
    end else begin
      deltas_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state175) | (1'b1 == ap_CS_fsm_state115) | (1'b1 == ap_CS_fsm_state179) | (1'b1 == ap_CS_fsm_state117) | (1'b1 == ap_CS_fsm_state67)) begin
      deltas_ce0 = 1'b1;
    end else begin
      deltas_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state175) | (1'b1 == ap_CS_fsm_state115)) begin
      deltas_d0 = reg_596;
    end else if(1'b1 == ap_CS_fsm_state67) begin
      deltas_d0 = 64'd0;
    end else begin
      deltas_d0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state175) | (1'b1 == ap_CS_fsm_state115) | (icmp_ln111_fu_1148_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state67)) begin
      deltas_we0 = 1'b1;
    end else begin
      deltas_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state70) begin
      grp_fu_559_opcode = 2'd1;
    end else if((1'b1 == ap_CS_fsm_state196) | (1'b1 == ap_CS_fsm_state191) | (1'b1 == ap_CS_fsm_state143) | (1'b1 == ap_CS_fsm_state124) | (1'b1 == ap_CS_fsm_state83) | (1'b1 == ap_CS_fsm_state38) | (1'b1 == ap_CS_fsm_state20)) begin
      grp_fu_559_opcode = 2'd0;
    end else begin
      grp_fu_559_opcode = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state196) begin
      grp_fu_559_p0 = reg_609;
    end else if(1'b1 == ap_CS_fsm_state191) begin
      grp_fu_559_p0 = reg_590;
    end else if(1'b1 == ap_CS_fsm_state124) begin
      grp_fu_559_p0 = error_0_i_i_0_reg_514;
    end else if(1'b1 == ap_CS_fsm_state70) begin
      grp_fu_559_p0 = targets_load_reg_1790;
    end else if((1'b1 == ap_CS_fsm_state143) | (1'b1 == ap_CS_fsm_state83) | (1'b1 == ap_CS_fsm_state38)) begin
      grp_fu_559_p0 = reg_604;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      grp_fu_559_p0 = x_assign_1_reg_447;
    end else begin
      grp_fu_559_p0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state70) begin
      grp_fu_559_p1 = reg_583;
    end else if((1'b1 == ap_CS_fsm_state143) | (1'b1 == ap_CS_fsm_state83) | (1'b1 == ap_CS_fsm_state38)) begin
      grp_fu_559_p1 = 64'd4607182418800017408;
    end else if((1'b1 == ap_CS_fsm_state196) | (1'b1 == ap_CS_fsm_state191) | (1'b1 == ap_CS_fsm_state124) | (1'b1 == ap_CS_fsm_state20)) begin
      grp_fu_559_p1 = reg_596;
    end else begin
      grp_fu_559_p1 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state191) begin
      grp_fu_566_p0 = changeMat_load_reg_1948;
    end else if(1'b1 == ap_CS_fsm_state186) begin
      grp_fu_566_p0 = reg_596;
    end else if((1'b1 == ap_CS_fsm_state181) | (1'b1 == ap_CS_fsm_state119)) begin
      grp_fu_566_p0 = reg_623;
    end else if((1'b1 == ap_CS_fsm_state170) | (1'b1 == ap_CS_fsm_state110)) begin
      grp_fu_566_p0 = reg_617;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      grp_fu_566_p0 = reg_583;
    end else begin
      grp_fu_566_p0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state191) begin
      grp_fu_566_p1 = 64'd4591870180066957722;
    end else if(1'b1 == ap_CS_fsm_state186) begin
      grp_fu_566_p1 = 64'd4602678819172646912;
    end else if(1'b1 == ap_CS_fsm_state181) begin
      grp_fu_566_p1 = reg_583;
    end else if(1'b1 == ap_CS_fsm_state170) begin
      grp_fu_566_p1 = error_0_i_i_0_reg_514;
    end else if(1'b1 == ap_CS_fsm_state110) begin
      grp_fu_566_p1 = reg_609;
    end else if((1'b1 == ap_CS_fsm_state119) | (1'b1 == ap_CS_fsm_state15)) begin
      grp_fu_566_p1 = reg_590;
    end else begin
      grp_fu_566_p1 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state88) begin
      grp_fu_573_p1 = temp_reg_1805;
    end else if((1'b1 == ap_CS_fsm_state148) | (1'b1 == ap_CS_fsm_state43)) begin
      grp_fu_573_p1 = reg_609;
    end else begin
      grp_fu_573_p1 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state130) begin
      grp_fu_578_p1 = bitcast_ln7_5_fu_1352_p1;
    end else if(1'b1 == ap_CS_fsm_state70) begin
      grp_fu_578_p1 = bitcast_ln7_1_fu_1225_p1;
    end else if(1'b1 == ap_CS_fsm_state25) begin
      grp_fu_578_p1 = bitcast_ln7_3_fu_1102_p1;
    end else begin
      grp_fu_578_p1 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      inputs_ce0 = 1'b1;
    end else begin
      inputs_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state68) begin
      targets_ce0 = 1'b1;
    end else begin
      targets_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state189) | (1'b1 == ap_CS_fsm_state201)) begin
      weights_address0 = weights_addr_2_reg_1933;
    end else if(1'b1 == ap_CS_fsm_state117) begin
      weights_address0 = zext_ln73_7_fu_1326_p1;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      weights_address0 = zext_ln21_5_fu_1087_p1;
    end else begin
      weights_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state189) | (1'b1 == ap_CS_fsm_state201) | (1'b1 == ap_CS_fsm_state117) | (1'b1 == ap_CS_fsm_state13)) begin
      weights_ce0 = 1'b1;
    end else begin
      weights_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state201) begin
      weights_we0 = 1'b1;
    end else begin
      weights_we0 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if((icmp_ln156_fu_628_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end
      end
      ap_ST_fsm_state3: begin
        if((icmp_ln157_fu_670_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state3)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end
      end
      ap_ST_fsm_state4: begin
        if((icmp_ln159_fu_726_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state4)) begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end
      end
      ap_ST_fsm_state5: begin
        if((icmp_ln165_fu_752_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state5)) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end
      end
      ap_ST_fsm_state6: begin
        if((icmp_ln167_fu_764_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state6)) begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end
      end
      ap_ST_fsm_state7: begin
        if((icmp_ln168_fu_776_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state7)) begin
          ap_NS_fsm = ap_ST_fsm_state9;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state8: begin
        if((icmp_ln169_fu_860_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state8)) begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state9: begin
        if((icmp_ln34_fu_886_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state9)) begin
          ap_NS_fsm = ap_ST_fsm_state11;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state10;
        end
      end
      ap_ST_fsm_state10: begin
        ap_NS_fsm = ap_ST_fsm_state9;
      end
      ap_ST_fsm_state11: begin
        if((icmp_ln39_fu_917_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state11)) begin
          ap_NS_fsm = ap_ST_fsm_state66;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state12;
        end
      end
      ap_ST_fsm_state12: begin
        if((icmp_ln18_fu_1001_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state12)) begin
          ap_NS_fsm = ap_ST_fsm_state11;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state13;
        end
      end
      ap_ST_fsm_state13: begin
        if((icmp_ln20_fu_1031_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state13)) begin
          ap_NS_fsm = ap_ST_fsm_state25;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state14;
        end
      end
      ap_ST_fsm_state14: begin
        begin
          if(working_key[0] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state184;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state15;
          end
        end
      end
      ap_ST_fsm_state15: begin
        begin
          if(working_key[1] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state16;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state77;
          end
        end
      end
      ap_ST_fsm_state16: begin
        begin
          if(working_key[2] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state97;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state17;
          end
        end
      end
      ap_ST_fsm_state17: begin
        begin
          if(working_key[3] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state116;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state18;
          end
        end
      end
      ap_ST_fsm_state18: begin
        begin
          if(working_key[4] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state19;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state127;
          end
        end
      end
      ap_ST_fsm_state19: begin
        begin
          if(working_key[5] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state80;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state20;
          end
        end
      end
      ap_ST_fsm_state20: begin
        begin
          if(working_key[6] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state120;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state21;
          end
        end
      end
      ap_ST_fsm_state21: begin
        begin
          if(working_key[7] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state22;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state181;
          end
        end
      end
      ap_ST_fsm_state22: begin
        begin
          if(working_key[8] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state23;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state119;
          end
        end
      end
      ap_ST_fsm_state23: begin
        begin
          if(working_key[9] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state24;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state154;
          end
        end
      end
      ap_ST_fsm_state24: begin
        begin
          if(working_key[10] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state114;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state13;
          end
        end
      end
      ap_ST_fsm_state25: begin
        begin
          if(working_key[11] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state132;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state26;
          end
        end
      end
      ap_ST_fsm_state26: begin
        begin
          if(working_key[12] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state27;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state140;
          end
        end
      end
      ap_ST_fsm_state27: begin
        begin
          if(working_key[13] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state33;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state28;
          end
        end
      end
      ap_ST_fsm_state28: begin
        begin
          if(working_key[14] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state29;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state57;
          end
        end
      end
      ap_ST_fsm_state29: begin
        begin
          if(working_key[15] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state30;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state33;
          end
        end
      end
      ap_ST_fsm_state30: begin
        begin
          if(working_key[16] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state28;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state31;
          end
        end
      end
      ap_ST_fsm_state31: begin
        begin
          if(working_key[17] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state131;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state32;
          end
        end
      end
      ap_ST_fsm_state32: begin
        begin
          if(working_key[18] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state33;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state133;
          end
        end
      end
      ap_ST_fsm_state33: begin
        begin
          if(working_key[19] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state34;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state185;
          end
        end
      end
      ap_ST_fsm_state34: begin
        begin
          if(working_key[20] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state35;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state60;
          end
        end
      end
      ap_ST_fsm_state35: begin
        begin
          if(working_key[21] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state140;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state36;
          end
        end
      end
      ap_ST_fsm_state36: begin
        begin
          if(working_key[22] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state37;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state47;
          end
        end
      end
      ap_ST_fsm_state37: begin
        begin
          if(working_key[23] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state42;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state38;
          end
        end
      end
      ap_ST_fsm_state38: begin
        begin
          if(working_key[24] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state149;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state39;
          end
        end
      end
      ap_ST_fsm_state39: begin
        begin
          if(working_key[25] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state200;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state40;
          end
        end
      end
      ap_ST_fsm_state40: begin
        begin
          if(working_key[26] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state41;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state73;
          end
        end
      end
      ap_ST_fsm_state41: begin
        begin
          if(working_key[27] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state129;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state42;
          end
        end
      end
      ap_ST_fsm_state42: begin
        begin
          if(working_key[28] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state29;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state43;
          end
        end
      end
      ap_ST_fsm_state43: begin
        begin
          if(working_key[29] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state154;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state44;
          end
        end
      end
      ap_ST_fsm_state44: begin
        begin
          if(working_key[30] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state45;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state165;
          end
        end
      end
      ap_ST_fsm_state45: begin
        begin
          if(working_key[31] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state46;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state101;
          end
        end
      end
      ap_ST_fsm_state46: begin
        begin
          if(working_key[32] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state60;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state47;
          end
        end
      end
      ap_ST_fsm_state47: begin
        begin
          if(working_key[33] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state48;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state170;
          end
        end
      end
      ap_ST_fsm_state48: begin
        begin
          if(working_key[34] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state49;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state154;
          end
        end
      end
      ap_ST_fsm_state49: begin
        begin
          if(working_key[35] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state174;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state50;
          end
        end
      end
      ap_ST_fsm_state50: begin
        begin
          if(working_key[36] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state89;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state51;
          end
        end
      end
      ap_ST_fsm_state51: begin
        begin
          if(working_key[37] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state105;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state52;
          end
        end
      end
      ap_ST_fsm_state52: begin
        begin
          if(working_key[38] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state53;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state73;
          end
        end
      end
      ap_ST_fsm_state53: begin
        begin
          if(working_key[39] == 1'b1) begin
            ap_NS_fsm = ap_ST_fsm_state54;
          end else begin
            ap_NS_fsm = ap_ST_fsm_state123;
          end
        end
      end
      ap_ST_fsm_state54: begin
        ap_NS_fsm = ap_ST_fsm_state55;
      end
      ap_ST_fsm_state55: begin
        ap_NS_fsm = ap_ST_fsm_state56;
      end
      ap_ST_fsm_state56: begin
        ap_NS_fsm = ap_ST_fsm_state57;
      end
      ap_ST_fsm_state57: begin
        ap_NS_fsm = ap_ST_fsm_state58;
      end
      ap_ST_fsm_state58: begin
        ap_NS_fsm = ap_ST_fsm_state59;
      end
      ap_ST_fsm_state59: begin
        ap_NS_fsm = ap_ST_fsm_state60;
      end
      ap_ST_fsm_state60: begin
        ap_NS_fsm = ap_ST_fsm_state61;
      end
      ap_ST_fsm_state61: begin
        ap_NS_fsm = ap_ST_fsm_state62;
      end
      ap_ST_fsm_state62: begin
        ap_NS_fsm = ap_ST_fsm_state63;
      end
      ap_ST_fsm_state63: begin
        ap_NS_fsm = ap_ST_fsm_state64;
      end
      ap_ST_fsm_state64: begin
        ap_NS_fsm = ap_ST_fsm_state65;
      end
      ap_ST_fsm_state65: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      ap_ST_fsm_state66: begin
        if((icmp_ln110_fu_1106_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state66)) begin
          ap_NS_fsm = ap_ST_fsm_state68;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state67;
        end
      end
      ap_ST_fsm_state67: begin
        if((icmp_ln111_fu_1148_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state67)) begin
          ap_NS_fsm = ap_ST_fsm_state66;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state67;
        end
      end
      ap_ST_fsm_state68: begin
        if((icmp_ln51_fu_1174_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state68)) begin
          ap_NS_fsm = ap_ST_fsm_state116;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state69;
        end
      end
      ap_ST_fsm_state69: begin
        ap_NS_fsm = ap_ST_fsm_state70;
      end
      ap_ST_fsm_state70: begin
        ap_NS_fsm = ap_ST_fsm_state71;
      end
      ap_ST_fsm_state71: begin
        ap_NS_fsm = ap_ST_fsm_state72;
      end
      ap_ST_fsm_state72: begin
        ap_NS_fsm = ap_ST_fsm_state73;
      end
      ap_ST_fsm_state73: begin
        ap_NS_fsm = ap_ST_fsm_state74;
      end
      ap_ST_fsm_state74: begin
        ap_NS_fsm = ap_ST_fsm_state75;
      end
      ap_ST_fsm_state75: begin
        ap_NS_fsm = ap_ST_fsm_state76;
      end
      ap_ST_fsm_state76: begin
        ap_NS_fsm = ap_ST_fsm_state77;
      end
      ap_ST_fsm_state77: begin
        ap_NS_fsm = ap_ST_fsm_state78;
      end
      ap_ST_fsm_state78: begin
        ap_NS_fsm = ap_ST_fsm_state79;
      end
      ap_ST_fsm_state79: begin
        ap_NS_fsm = ap_ST_fsm_state80;
      end
      ap_ST_fsm_state80: begin
        ap_NS_fsm = ap_ST_fsm_state81;
      end
      ap_ST_fsm_state81: begin
        ap_NS_fsm = ap_ST_fsm_state82;
      end
      ap_ST_fsm_state82: begin
        ap_NS_fsm = ap_ST_fsm_state83;
      end
      ap_ST_fsm_state83: begin
        ap_NS_fsm = ap_ST_fsm_state84;
      end
      ap_ST_fsm_state84: begin
        ap_NS_fsm = ap_ST_fsm_state85;
      end
      ap_ST_fsm_state85: begin
        ap_NS_fsm = ap_ST_fsm_state86;
      end
      ap_ST_fsm_state86: begin
        ap_NS_fsm = ap_ST_fsm_state87;
      end
      ap_ST_fsm_state87: begin
        ap_NS_fsm = ap_ST_fsm_state88;
      end
      ap_ST_fsm_state88: begin
        ap_NS_fsm = ap_ST_fsm_state89;
      end
      ap_ST_fsm_state89: begin
        ap_NS_fsm = ap_ST_fsm_state90;
      end
      ap_ST_fsm_state90: begin
        ap_NS_fsm = ap_ST_fsm_state91;
      end
      ap_ST_fsm_state91: begin
        ap_NS_fsm = ap_ST_fsm_state92;
      end
      ap_ST_fsm_state92: begin
        ap_NS_fsm = ap_ST_fsm_state93;
      end
      ap_ST_fsm_state93: begin
        ap_NS_fsm = ap_ST_fsm_state94;
      end
      ap_ST_fsm_state94: begin
        ap_NS_fsm = ap_ST_fsm_state95;
      end
      ap_ST_fsm_state95: begin
        ap_NS_fsm = ap_ST_fsm_state96;
      end
      ap_ST_fsm_state96: begin
        ap_NS_fsm = ap_ST_fsm_state97;
      end
      ap_ST_fsm_state97: begin
        ap_NS_fsm = ap_ST_fsm_state98;
      end
      ap_ST_fsm_state98: begin
        ap_NS_fsm = ap_ST_fsm_state99;
      end
      ap_ST_fsm_state99: begin
        ap_NS_fsm = ap_ST_fsm_state100;
      end
      ap_ST_fsm_state100: begin
        ap_NS_fsm = ap_ST_fsm_state101;
      end
      ap_ST_fsm_state101: begin
        ap_NS_fsm = ap_ST_fsm_state102;
      end
      ap_ST_fsm_state102: begin
        ap_NS_fsm = ap_ST_fsm_state103;
      end
      ap_ST_fsm_state103: begin
        ap_NS_fsm = ap_ST_fsm_state104;
      end
      ap_ST_fsm_state104: begin
        ap_NS_fsm = ap_ST_fsm_state105;
      end
      ap_ST_fsm_state105: begin
        ap_NS_fsm = ap_ST_fsm_state106;
      end
      ap_ST_fsm_state106: begin
        ap_NS_fsm = ap_ST_fsm_state107;
      end
      ap_ST_fsm_state107: begin
        ap_NS_fsm = ap_ST_fsm_state108;
      end
      ap_ST_fsm_state108: begin
        ap_NS_fsm = ap_ST_fsm_state109;
      end
      ap_ST_fsm_state109: begin
        ap_NS_fsm = ap_ST_fsm_state110;
      end
      ap_ST_fsm_state110: begin
        ap_NS_fsm = ap_ST_fsm_state111;
      end
      ap_ST_fsm_state111: begin
        ap_NS_fsm = ap_ST_fsm_state112;
      end
      ap_ST_fsm_state112: begin
        ap_NS_fsm = ap_ST_fsm_state113;
      end
      ap_ST_fsm_state113: begin
        ap_NS_fsm = ap_ST_fsm_state114;
      end
      ap_ST_fsm_state114: begin
        ap_NS_fsm = ap_ST_fsm_state115;
      end
      ap_ST_fsm_state115: begin
        ap_NS_fsm = ap_ST_fsm_state68;
      end
      ap_ST_fsm_state116: begin
        if((icmp_ln70_fu_1239_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state116)) begin
          ap_NS_fsm = ap_ST_fsm_state176;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state117;
        end
      end
      ap_ST_fsm_state117: begin
        if((icmp_ln72_fu_1301_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state117)) begin
          ap_NS_fsm = ap_ST_fsm_state129;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state118;
        end
      end
      ap_ST_fsm_state118: begin
        ap_NS_fsm = ap_ST_fsm_state119;
      end
      ap_ST_fsm_state119: begin
        ap_NS_fsm = ap_ST_fsm_state120;
      end
      ap_ST_fsm_state120: begin
        ap_NS_fsm = ap_ST_fsm_state121;
      end
      ap_ST_fsm_state121: begin
        ap_NS_fsm = ap_ST_fsm_state122;
      end
      ap_ST_fsm_state122: begin
        ap_NS_fsm = ap_ST_fsm_state123;
      end
      ap_ST_fsm_state123: begin
        ap_NS_fsm = ap_ST_fsm_state124;
      end
      ap_ST_fsm_state124: begin
        ap_NS_fsm = ap_ST_fsm_state125;
      end
      ap_ST_fsm_state125: begin
        ap_NS_fsm = ap_ST_fsm_state126;
      end
      ap_ST_fsm_state126: begin
        ap_NS_fsm = ap_ST_fsm_state127;
      end
      ap_ST_fsm_state127: begin
        ap_NS_fsm = ap_ST_fsm_state128;
      end
      ap_ST_fsm_state128: begin
        ap_NS_fsm = ap_ST_fsm_state117;
      end
      ap_ST_fsm_state129: begin
        ap_NS_fsm = ap_ST_fsm_state130;
      end
      ap_ST_fsm_state130: begin
        ap_NS_fsm = ap_ST_fsm_state131;
      end
      ap_ST_fsm_state131: begin
        ap_NS_fsm = ap_ST_fsm_state132;
      end
      ap_ST_fsm_state132: begin
        ap_NS_fsm = ap_ST_fsm_state133;
      end
      ap_ST_fsm_state133: begin
        ap_NS_fsm = ap_ST_fsm_state134;
      end
      ap_ST_fsm_state134: begin
        ap_NS_fsm = ap_ST_fsm_state135;
      end
      ap_ST_fsm_state135: begin
        ap_NS_fsm = ap_ST_fsm_state136;
      end
      ap_ST_fsm_state136: begin
        ap_NS_fsm = ap_ST_fsm_state137;
      end
      ap_ST_fsm_state137: begin
        ap_NS_fsm = ap_ST_fsm_state138;
      end
      ap_ST_fsm_state138: begin
        ap_NS_fsm = ap_ST_fsm_state139;
      end
      ap_ST_fsm_state139: begin
        ap_NS_fsm = ap_ST_fsm_state140;
      end
      ap_ST_fsm_state140: begin
        ap_NS_fsm = ap_ST_fsm_state141;
      end
      ap_ST_fsm_state141: begin
        ap_NS_fsm = ap_ST_fsm_state142;
      end
      ap_ST_fsm_state142: begin
        ap_NS_fsm = ap_ST_fsm_state143;
      end
      ap_ST_fsm_state143: begin
        ap_NS_fsm = ap_ST_fsm_state144;
      end
      ap_ST_fsm_state144: begin
        ap_NS_fsm = ap_ST_fsm_state145;
      end
      ap_ST_fsm_state145: begin
        ap_NS_fsm = ap_ST_fsm_state146;
      end
      ap_ST_fsm_state146: begin
        ap_NS_fsm = ap_ST_fsm_state147;
      end
      ap_ST_fsm_state147: begin
        ap_NS_fsm = ap_ST_fsm_state148;
      end
      ap_ST_fsm_state148: begin
        ap_NS_fsm = ap_ST_fsm_state149;
      end
      ap_ST_fsm_state149: begin
        ap_NS_fsm = ap_ST_fsm_state150;
      end
      ap_ST_fsm_state150: begin
        ap_NS_fsm = ap_ST_fsm_state151;
      end
      ap_ST_fsm_state151: begin
        ap_NS_fsm = ap_ST_fsm_state152;
      end
      ap_ST_fsm_state152: begin
        ap_NS_fsm = ap_ST_fsm_state153;
      end
      ap_ST_fsm_state153: begin
        ap_NS_fsm = ap_ST_fsm_state154;
      end
      ap_ST_fsm_state154: begin
        ap_NS_fsm = ap_ST_fsm_state155;
      end
      ap_ST_fsm_state155: begin
        ap_NS_fsm = ap_ST_fsm_state156;
      end
      ap_ST_fsm_state156: begin
        ap_NS_fsm = ap_ST_fsm_state157;
      end
      ap_ST_fsm_state157: begin
        ap_NS_fsm = ap_ST_fsm_state158;
      end
      ap_ST_fsm_state158: begin
        ap_NS_fsm = ap_ST_fsm_state159;
      end
      ap_ST_fsm_state159: begin
        ap_NS_fsm = ap_ST_fsm_state160;
      end
      ap_ST_fsm_state160: begin
        ap_NS_fsm = ap_ST_fsm_state161;
      end
      ap_ST_fsm_state161: begin
        ap_NS_fsm = ap_ST_fsm_state162;
      end
      ap_ST_fsm_state162: begin
        ap_NS_fsm = ap_ST_fsm_state163;
      end
      ap_ST_fsm_state163: begin
        ap_NS_fsm = ap_ST_fsm_state164;
      end
      ap_ST_fsm_state164: begin
        ap_NS_fsm = ap_ST_fsm_state165;
      end
      ap_ST_fsm_state165: begin
        ap_NS_fsm = ap_ST_fsm_state166;
      end
      ap_ST_fsm_state166: begin
        ap_NS_fsm = ap_ST_fsm_state167;
      end
      ap_ST_fsm_state167: begin
        ap_NS_fsm = ap_ST_fsm_state168;
      end
      ap_ST_fsm_state168: begin
        ap_NS_fsm = ap_ST_fsm_state169;
      end
      ap_ST_fsm_state169: begin
        ap_NS_fsm = ap_ST_fsm_state170;
      end
      ap_ST_fsm_state170: begin
        ap_NS_fsm = ap_ST_fsm_state171;
      end
      ap_ST_fsm_state171: begin
        ap_NS_fsm = ap_ST_fsm_state172;
      end
      ap_ST_fsm_state172: begin
        ap_NS_fsm = ap_ST_fsm_state173;
      end
      ap_ST_fsm_state173: begin
        ap_NS_fsm = ap_ST_fsm_state174;
      end
      ap_ST_fsm_state174: begin
        ap_NS_fsm = ap_ST_fsm_state175;
      end
      ap_ST_fsm_state175: begin
        ap_NS_fsm = ap_ST_fsm_state116;
      end
      ap_ST_fsm_state176: begin
        if((icmp_ln123_fu_1356_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state176)) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state177;
        end
      end
      ap_ST_fsm_state177: begin
        if((icmp_ln87_fu_1442_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state177)) begin
          ap_NS_fsm = ap_ST_fsm_state176;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state178;
        end
      end
      ap_ST_fsm_state178: begin
        ap_NS_fsm = ap_ST_fsm_state179;
      end
      ap_ST_fsm_state179: begin
        if((icmp_ln88_fu_1524_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state179)) begin
          ap_NS_fsm = ap_ST_fsm_state177;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state180;
        end
      end
      ap_ST_fsm_state180: begin
        ap_NS_fsm = ap_ST_fsm_state181;
      end
      ap_ST_fsm_state181: begin
        ap_NS_fsm = ap_ST_fsm_state182;
      end
      ap_ST_fsm_state182: begin
        ap_NS_fsm = ap_ST_fsm_state183;
      end
      ap_ST_fsm_state183: begin
        ap_NS_fsm = ap_ST_fsm_state184;
      end
      ap_ST_fsm_state184: begin
        ap_NS_fsm = ap_ST_fsm_state185;
      end
      ap_ST_fsm_state185: begin
        ap_NS_fsm = ap_ST_fsm_state186;
      end
      ap_ST_fsm_state186: begin
        ap_NS_fsm = ap_ST_fsm_state187;
      end
      ap_ST_fsm_state187: begin
        ap_NS_fsm = ap_ST_fsm_state188;
      end
      ap_ST_fsm_state188: begin
        ap_NS_fsm = ap_ST_fsm_state189;
      end
      ap_ST_fsm_state189: begin
        ap_NS_fsm = ap_ST_fsm_state190;
      end
      ap_ST_fsm_state190: begin
        ap_NS_fsm = ap_ST_fsm_state191;
      end
      ap_ST_fsm_state191: begin
        ap_NS_fsm = ap_ST_fsm_state192;
      end
      ap_ST_fsm_state192: begin
        ap_NS_fsm = ap_ST_fsm_state193;
      end
      ap_ST_fsm_state193: begin
        ap_NS_fsm = ap_ST_fsm_state194;
      end
      ap_ST_fsm_state194: begin
        ap_NS_fsm = ap_ST_fsm_state195;
      end
      ap_ST_fsm_state195: begin
        ap_NS_fsm = ap_ST_fsm_state196;
      end
      ap_ST_fsm_state196: begin
        ap_NS_fsm = ap_ST_fsm_state197;
      end
      ap_ST_fsm_state197: begin
        ap_NS_fsm = ap_ST_fsm_state198;
      end
      ap_ST_fsm_state198: begin
        ap_NS_fsm = ap_ST_fsm_state199;
      end
      ap_ST_fsm_state199: begin
        ap_NS_fsm = ap_ST_fsm_state200;
      end
      ap_ST_fsm_state200: begin
        ap_NS_fsm = ap_ST_fsm_state201;
      end
      ap_ST_fsm_state201: begin
        ap_NS_fsm = ap_ST_fsm_state179;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign add_ln112_1_fu_1164_p2 = add_ln112_reg_1754 + zext_ln112_2_fu_1160_p1;
  assign add_ln112_fu_1142_p2 = zext_ln112_1_fu_1138_p1 + zext_ln112_fu_1126_p1;
  assign add_ln160_1_fu_686_p2 = zext_ln160_2_fu_682_p1 + add_ln160_reg_1586;
  assign add_ln160_2_fu_720_p2 = zext_ln160_4_fu_704_p1 + zext_ln160_5_fu_716_p1;
  assign add_ln160_3_fu_742_p2 = add_ln160_2_reg_1599 + zext_ln160_6_fu_738_p1;
  assign add_ln160_fu_664_p2 = zext_ln160_1_fu_660_p1 + zext_ln160_fu_648_p1;
  assign add_ln170_1_fu_876_p2 = add_ln170_reg_1636 + zext_ln170_2_fu_872_p1;
  assign add_ln170_fu_812_p2 = zext_ln170_1_fu_808_p1 + zext_ln170_fu_796_p1;
  assign add_ln21_1_fu_1046_p2 = zext_ln21_2_fu_1042_p1 + add_ln21_reg_1680;
  assign add_ln21_2_fu_1076_p2 = p_shl_cast_fu_1056_p3 + zext_ln21_4_fu_1072_p1;
  assign add_ln21_3_fu_1082_p2 = zext_ln23_2_reg_1703 + add_ln21_2_fu_1076_p2;
  assign add_ln21_fu_953_p2 = zext_ln21_fu_937_p1 + zext_ln21_1_fu_949_p1;
  assign add_ln23_1_fu_1021_p2 = add_ln23_reg_1690 + zext_ln23_3_fu_1017_p1;
  assign add_ln23_fu_995_p2 = zext_ln23_fu_979_p1 + zext_ln23_1_fu_991_p1;
  assign add_ln35_fu_902_p2 = zext_ln52_reg_1641 + zext_ln35_1_fu_898_p1;
  assign add_ln52_1_fu_1194_p2 = add_ln52_reg_1646 + zext_ln52_4_fu_1190_p1;
  assign add_ln52_2_fu_1204_p2 = $signed(zext_ln52_3_fu_1186_p1) + $signed(5'd20);
  assign add_ln52_fu_854_p2 = zext_ln52_2_fu_850_p1 + zext_ln52_1_fu_838_p1;
  assign add_ln53_fu_1229_p2 = zext_ln52_3_reg_1775 + 5'd10;
  assign add_ln70_fu_1245_p2 = jj_0_i_i21_0_reg_492 + 4'd1;
  assign add_ln72_fu_1307_p2 = kk_0_i_i_0_reg_503 + 4'd1;
  assign add_ln73_1_fu_1295_p2 = zext_ln73_3_fu_1279_p1 + zext_ln73_4_fu_1291_p1;
  assign add_ln73_2_fu_1321_p2 = add_ln73_1_reg_1818 + zext_ln73_6_fu_1317_p1;
  assign add_ln73_3_fu_1331_p2 = zext_ln73_5_fu_1313_p1 + 5'd10;
  assign add_ln73_fu_1260_p2 = zext_ln73_1_fu_1256_p1 + 5'd10;
  assign add_ln89_fu_1558_p2 = add_ln90_reg_1874 + zext_ln90_10_fu_1540_p1;
  assign add_ln90_1_fu_1422_p2 = zext_ln90_3_fu_1418_p1 + zext_ln90_2_fu_1406_p1;
  assign add_ln90_2_fu_1457_p2 = zext_ln90_4_fu_1453_p1 + add_ln90_reg_1874;
  assign add_ln90_3_fu_1490_p2 = p_shl6_cast_fu_1472_p3 + zext_ln90_6_fu_1486_p1;
  assign add_ln90_4_fu_1467_p2 = zext_ln90_4_fu_1453_p1 + add_ln90_1_reg_1880;
  assign add_ln90_5_fu_1518_p2 = zext_ln90_7_fu_1503_p1 + zext_ln90_8_fu_1514_p1;
  assign add_ln90_6_fu_1548_p2 = add_ln90_3_reg_1915 + zext_ln90_11_fu_1544_p1;
  assign add_ln90_7_fu_1568_p2 = add_ln90_5_reg_1920 + zext_ln90_9_fu_1536_p1;
  assign add_ln90_fu_1392_p2 = zext_ln90_1_fu_1388_p1 + zext_ln90_fu_1376_p1;
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state109 = ap_CS_fsm[32'd108];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state110 = ap_CS_fsm[32'd109];
  assign ap_CS_fsm_state114 = ap_CS_fsm[32'd113];
  assign ap_CS_fsm_state115 = ap_CS_fsm[32'd114];
  assign ap_CS_fsm_state116 = ap_CS_fsm[32'd115];
  assign ap_CS_fsm_state117 = ap_CS_fsm[32'd116];
  assign ap_CS_fsm_state118 = ap_CS_fsm[32'd117];
  assign ap_CS_fsm_state119 = ap_CS_fsm[32'd118];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state123 = ap_CS_fsm[32'd122];
  assign ap_CS_fsm_state124 = ap_CS_fsm[32'd123];
  assign ap_CS_fsm_state128 = ap_CS_fsm[32'd127];
  assign ap_CS_fsm_state129 = ap_CS_fsm[32'd128];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state130 = ap_CS_fsm[32'd129];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state142 = ap_CS_fsm[32'd141];
  assign ap_CS_fsm_state143 = ap_CS_fsm[32'd142];
  assign ap_CS_fsm_state147 = ap_CS_fsm[32'd146];
  assign ap_CS_fsm_state148 = ap_CS_fsm[32'd147];
  assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];
  assign ap_CS_fsm_state169 = ap_CS_fsm[32'd168];
  assign ap_CS_fsm_state170 = ap_CS_fsm[32'd169];
  assign ap_CS_fsm_state174 = ap_CS_fsm[32'd173];
  assign ap_CS_fsm_state175 = ap_CS_fsm[32'd174];
  assign ap_CS_fsm_state176 = ap_CS_fsm[32'd175];
  assign ap_CS_fsm_state177 = ap_CS_fsm[32'd176];
  assign ap_CS_fsm_state178 = ap_CS_fsm[32'd177];
  assign ap_CS_fsm_state179 = ap_CS_fsm[32'd178];
  assign ap_CS_fsm_state180 = ap_CS_fsm[32'd179];
  assign ap_CS_fsm_state181 = ap_CS_fsm[32'd180];
  assign ap_CS_fsm_state185 = ap_CS_fsm[32'd184];
  assign ap_CS_fsm_state186 = ap_CS_fsm[32'd185];
  assign ap_CS_fsm_state187 = ap_CS_fsm[32'd186];
  assign ap_CS_fsm_state189 = ap_CS_fsm[32'd188];
  assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];
  assign ap_CS_fsm_state190 = ap_CS_fsm[32'd189];
  assign ap_CS_fsm_state191 = ap_CS_fsm[32'd190];
  assign ap_CS_fsm_state195 = ap_CS_fsm[32'd194];
  assign ap_CS_fsm_state196 = ap_CS_fsm[32'd195];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];
  assign ap_CS_fsm_state200 = ap_CS_fsm[32'd199];
  assign ap_CS_fsm_state201 = ap_CS_fsm[32'd200];
  assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];
  assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state37 = ap_CS_fsm[32'd36];
  assign ap_CS_fsm_state38 = ap_CS_fsm[32'd37];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state42 = ap_CS_fsm[32'd41];
  assign ap_CS_fsm_state43 = ap_CS_fsm[32'd42];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state64 = ap_CS_fsm[32'd63];
  assign ap_CS_fsm_state65 = ap_CS_fsm[32'd64];
  assign ap_CS_fsm_state66 = ap_CS_fsm[32'd65];
  assign ap_CS_fsm_state67 = ap_CS_fsm[32'd66];
  assign ap_CS_fsm_state68 = ap_CS_fsm[32'd67];
  assign ap_CS_fsm_state69 = ap_CS_fsm[32'd68];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state70 = ap_CS_fsm[32'd69];
  assign ap_CS_fsm_state74 = ap_CS_fsm[32'd73];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state82 = ap_CS_fsm[32'd81];
  assign ap_CS_fsm_state83 = ap_CS_fsm[32'd82];
  assign ap_CS_fsm_state87 = ap_CS_fsm[32'd86];
  assign ap_CS_fsm_state88 = ap_CS_fsm[32'd87];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign bitcast_ln7_1_fu_1225_p1 = xor_ln7_reg_1795;
  assign bitcast_ln7_2_fu_1092_p1 = x_assign_1_reg_447;
  assign bitcast_ln7_3_fu_1102_p1 = xor_ln7_1_reg_1731;
  assign bitcast_ln7_4_fu_1342_p1 = activations_q0;
  assign bitcast_ln7_5_fu_1352_p1 = xor_ln7_2_reg_1856;
  assign bitcast_ln7_fu_1215_p1 = activations_q0;
  assign cols_2_fu_782_p2 = cols_1_reg_380 + 2'd1;
  assign cols_fu_732_p2 = cols_0_reg_346 + 4'd1;
  assign ee_2_fu_758_p2 = ee_1_reg_357 + 7'd1;
  assign ee_fu_634_p2 = ee_0_reg_324 + 2'd1;
  assign i_1_fu_923_p2 = i_1_i_reg_414 + 2'd1;
  assign i_2_fu_1180_p2 = i_0_i_i_reg_481 + 4'd1;
  assign i_3_fu_1112_p2 = i_0_i13_reg_459 + 2'd1;
  assign i_fu_892_p2 = i_0_i_reg_402 + 3'd1;
  assign icmp_ln110_fu_1106_p2 = (i_0_i13_reg_459 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln111_fu_1148_p2 = (j_0_i_reg_470 == 4'd10)? 1'b1 : 1'b0;
  assign icmp_ln123_fu_1356_p2 = (level_assign_reg_526 == 2'd0)? 1'b1 : 1'b0;
  assign icmp_ln156_fu_628_p2 = (ee_0_reg_324 == 2'd3)? 1'b1 : 1'b0;
  assign icmp_ln157_fu_670_p2 = (rows_0_reg_335 == 4'd10)? 1'b1 : 1'b0;
  assign icmp_ln159_fu_726_p2 = (cols_0_reg_346 == 4'd10)? 1'b1 : 1'b0;
  assign icmp_ln165_fu_752_p2 = (ee_1_reg_357 == 7'd100)? 1'b1 : 1'b0;
  assign icmp_ln167_fu_764_p2 = (jj_0_reg_368 == 7'd100)? 1'b1 : 1'b0;
  assign icmp_ln168_fu_776_p2 = (cols_1_reg_380 == 2'd3)? 1'b1 : 1'b0;
  assign icmp_ln169_fu_860_p2 = (rows_1_reg_391 == 4'd10)? 1'b1 : 1'b0;
  assign icmp_ln18_fu_1001_p2 = (ii_0_i_i_reg_425 == 4'd10)? 1'b1 : 1'b0;
  assign icmp_ln20_fu_1031_p2 = (jj_0_i_i_reg_436 < select_ln40_reg_1685)? 1'b1 : 1'b0;
  assign icmp_ln34_fu_886_p2 = (i_0_i_reg_402 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln39_fu_917_p2 = (i_1_i_reg_414 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln51_fu_1174_p2 = (i_0_i_i_reg_481 == 4'd10)? 1'b1 : 1'b0;
  assign icmp_ln70_fu_1239_p2 = (jj_0_i_i21_0_reg_492 == 4'd10)? 1'b1 : 1'b0;
  assign icmp_ln72_fu_1301_p2 = (kk_0_i_i_0_reg_503 == 4'd10)? 1'b1 : 1'b0;
  assign icmp_ln87_1_fu_1428_p2 = (level_assign_reg_526 == 2'd1)? 1'b1 : 1'b0;
  assign icmp_ln87_fu_1442_p2 = (ii_0_i_i25_reg_537 < select_ln87_reg_1885)? 1'b1 : 1'b0;
  assign icmp_ln88_fu_1524_p2 = (jj_0_i10_i_reg_548 == 4'd10)? 1'b1 : 1'b0;
  assign ii_1_fu_1447_p2 = ii_0_i_i25_reg_537 + 4'd1;
  assign ii_fu_1007_p2 = ii_0_i_i_reg_425 + 4'd1;
  assign inputs_address0 = zext_ln35_2_fu_907_p1;
  assign j_2_fu_1362_p2 = $signed(level_assign_reg_526) + $signed(2'd3);
  assign j_fu_1154_p2 = j_0_i_reg_470 + 4'd1;
  assign jj_1_fu_770_p2 = jj_0_reg_368 + 7'd1;
  assign jj_2_fu_1530_p2 = jj_0_i10_i_reg_548 + 4'd1;
  assign jj_fu_1036_p2 = jj_0_i_i_reg_436 + 4'd1;
  assign p_shl6_cast_fu_1472_p3 = { { add_ln90_2_reg_1898 }, { 3'd0 } };
  assign p_shl_cast_fu_1056_p3 = { { add_ln21_1_fu_1046_p2 }, { 3'd0 } };
  assign rows_2_fu_866_p2 = rows_1_reg_391 + 4'd1;
  assign rows_fu_676_p2 = rows_0_reg_335 + 4'd1;
  assign select_ln40_fu_963_p3 = (trunc_ln40_fu_959_p1[0:0] === 1'b1)? 4'd10 : 4'd4;
  assign select_ln87_fu_1434_p3 = (icmp_ln87_1_fu_1428_p2[0:0] === 1'b1)? 4'd4 : 4'd10;
  assign targets_address0 = zext_ln52_5_fu_1199_p1;
  assign tmp_19_fu_652_p3 = { { ee_0_reg_324 }, { 1'd0 } };
  assign tmp_20_fu_696_p3 = { { add_ln160_1_fu_686_p2 }, { 3'd0 } };
  assign tmp_21_fu_708_p3 = { { add_ln160_1_fu_686_p2 }, { 1'd0 } };
  assign tmp_22_fu_818_p3 = { { jj_0_reg_368 }, { 2'd0 } };
  assign tmp_23_fu_830_p3 = { { jj_0_reg_368 }, { 3'd0 } };
  assign tmp_24_fu_842_p3 = { { jj_0_reg_368 }, { 1'd0 } };
  assign tmp_25_fu_788_p3 = { { cols_1_reg_380 }, { 3'd0 } };
  assign tmp_26_fu_800_p3 = { { cols_1_reg_380 }, { 1'd0 } };
  assign tmp_27_fu_929_p3 = { { i_1_i_reg_414 }, { 3'd0 } };
  assign tmp_28_fu_941_p3 = { { i_1_i_reg_414 }, { 1'd0 } };
  assign tmp_29_fu_971_p3 = { { i_1_fu_923_p2 }, { 3'd0 } };
  assign tmp_30_fu_983_p3 = { { i_1_fu_923_p2 }, { 1'd0 } };
  assign tmp_31_fu_1118_p3 = { { i_0_i13_reg_459 }, { 3'd0 } };
  assign tmp_32_fu_1130_p3 = { { i_0_i13_reg_459 }, { 1'd0 } };
  assign tmp_33_fu_1064_p3 = { { add_ln21_1_fu_1046_p2 }, { 1'd0 } };
  assign tmp_34_fu_1271_p3 = { { add_ln73_fu_1260_p2 }, { 3'd0 } };
  assign tmp_35_fu_1283_p3 = { { add_ln73_fu_1260_p2 }, { 1'd0 } };
  assign tmp_36_fu_1368_p3 = { { j_2_fu_1362_p2 }, { 3'd0 } };
  assign tmp_37_fu_1380_p3 = { { j_2_fu_1362_p2 }, { 1'd0 } };
  assign tmp_38_fu_1398_p3 = { { level_assign_reg_526 }, { 3'd0 } };
  assign tmp_39_fu_1410_p3 = { { level_assign_reg_526 }, { 1'd0 } };
  assign tmp_40_fu_1479_p3 = { { add_ln90_2_reg_1898 }, { 1'd0 } };
  assign tmp_41_fu_1496_p3 = { { add_ln90_4_reg_1904 }, { 3'd0 } };
  assign tmp_42_fu_1507_p3 = { { add_ln90_4_reg_1904 }, { 1'd0 } };
  assign tmp_fu_640_p3 = { { ee_0_reg_324 }, { 3'd0 } };
  assign trunc_ln40_fu_959_p1 = i_1_i_reg_414[0:0];
  assign weights_d0 = reg_609;
  assign xor_ln7_1_fu_1096_p2 = bitcast_ln7_2_fu_1092_p1 ^ 64'd9223372036854775808;
  assign xor_ln7_2_fu_1346_p2 = bitcast_ln7_4_fu_1342_p1 ^ 64'd9223372036854775808;
  assign xor_ln7_fu_1219_p2 = bitcast_ln7_fu_1215_p1 ^ 64'd9223372036854775808;
  assign zext_ln112_1_fu_1138_p1 = tmp_32_fu_1130_p3;
  assign zext_ln112_2_fu_1160_p1 = j_0_i_reg_470;
  assign zext_ln112_3_fu_1169_p1 = add_ln112_1_fu_1164_p2;
  assign zext_ln112_fu_1126_p1 = tmp_31_fu_1118_p3;
  assign zext_ln160_1_fu_660_p1 = tmp_19_fu_652_p3;
  assign zext_ln160_2_fu_682_p1 = rows_0_reg_335;
  assign zext_ln160_3_fu_691_p1 = add_ln160_1_fu_686_p2;
  assign zext_ln160_4_fu_704_p1 = tmp_20_fu_696_p3;
  assign zext_ln160_5_fu_716_p1 = tmp_21_fu_708_p3;
  assign zext_ln160_6_fu_738_p1 = cols_0_reg_346;
  assign zext_ln160_7_fu_747_p1 = add_ln160_3_fu_742_p2;
  assign zext_ln160_fu_648_p1 = tmp_fu_640_p3;
  assign zext_ln170_1_fu_808_p1 = tmp_26_fu_800_p3;
  assign zext_ln170_2_fu_872_p1 = rows_1_reg_391;
  assign zext_ln170_3_fu_881_p1 = add_ln170_1_fu_876_p2;
  assign zext_ln170_fu_796_p1 = tmp_25_fu_788_p3;
  assign zext_ln21_1_fu_949_p1 = tmp_28_fu_941_p3;
  assign zext_ln21_2_fu_1042_p1 = jj_0_i_i_reg_436;
  assign zext_ln21_3_fu_1051_p1 = add_ln21_1_fu_1046_p2;
  assign zext_ln21_4_fu_1072_p1 = tmp_33_fu_1064_p3;
  assign zext_ln21_5_fu_1087_p1 = add_ln21_3_fu_1082_p2;
  assign zext_ln21_fu_937_p1 = tmp_27_fu_929_p3;
  assign zext_ln23_1_fu_991_p1 = tmp_30_fu_983_p3;
  assign zext_ln23_2_fu_1013_p1 = ii_0_i_i_reg_425;
  assign zext_ln23_3_fu_1017_p1 = ii_0_i_i_reg_425;
  assign zext_ln23_4_fu_1026_p1 = add_ln23_1_fu_1021_p2;
  assign zext_ln23_fu_979_p1 = tmp_29_fu_971_p3;
  assign zext_ln35_1_fu_898_p1 = i_0_i_reg_402;
  assign zext_ln35_2_fu_907_p1 = add_ln35_fu_902_p2;
  assign zext_ln35_fu_912_p1 = i_0_i_reg_402;
  assign zext_ln52_1_fu_838_p1 = tmp_23_fu_830_p3;
  assign zext_ln52_2_fu_850_p1 = tmp_24_fu_842_p3;
  assign zext_ln52_3_fu_1186_p1 = i_0_i_i_reg_481;
  assign zext_ln52_4_fu_1190_p1 = i_0_i_i_reg_481;
  assign zext_ln52_5_fu_1199_p1 = add_ln52_1_fu_1194_p2;
  assign zext_ln52_6_fu_1210_p1 = add_ln52_2_fu_1204_p2;
  assign zext_ln52_fu_826_p1 = tmp_22_fu_818_p3;
  assign zext_ln53_fu_1234_p1 = add_ln53_fu_1229_p2;
  assign zext_ln73_1_fu_1256_p1 = jj_0_i_i21_0_reg_492;
  assign zext_ln73_2_fu_1266_p1 = add_ln73_fu_1260_p2;
  assign zext_ln73_3_fu_1279_p1 = tmp_34_fu_1271_p3;
  assign zext_ln73_4_fu_1291_p1 = tmp_35_fu_1283_p3;
  assign zext_ln73_5_fu_1313_p1 = kk_0_i_i_0_reg_503;
  assign zext_ln73_6_fu_1317_p1 = kk_0_i_i_0_reg_503;
  assign zext_ln73_7_fu_1326_p1 = add_ln73_2_fu_1321_p2;
  assign zext_ln73_8_fu_1337_p1 = add_ln73_3_fu_1331_p2;
  assign zext_ln73_fu_1251_p1 = jj_0_i_i21_0_reg_492;
  assign zext_ln89_fu_1563_p1 = add_ln89_fu_1558_p2;
  assign zext_ln90_10_fu_1540_p1 = jj_0_i10_i_reg_548;
  assign zext_ln90_11_fu_1544_p1 = jj_0_i10_i_reg_548;
  assign zext_ln90_12_fu_1553_p1 = add_ln90_6_fu_1548_p2;
  assign zext_ln90_13_fu_1573_p1 = add_ln90_7_fu_1568_p2;
  assign zext_ln90_1_fu_1388_p1 = tmp_37_fu_1380_p3;
  assign zext_ln90_2_fu_1406_p1 = tmp_38_fu_1398_p3;
  assign zext_ln90_3_fu_1418_p1 = tmp_39_fu_1410_p3;
  assign zext_ln90_4_fu_1453_p1 = ii_0_i_i25_reg_537;
  assign zext_ln90_5_fu_1462_p1 = add_ln90_2_fu_1457_p2;
  assign zext_ln90_6_fu_1486_p1 = tmp_40_fu_1479_p3;
  assign zext_ln90_7_fu_1503_p1 = tmp_41_fu_1496_p3;
  assign zext_ln90_8_fu_1514_p1 = tmp_42_fu_1507_p3;
  assign zext_ln90_9_fu_1536_p1 = jj_0_i10_i_reg_548;
  assign zext_ln90_fu_1376_p1 = tmp_36_fu_1368_p3;

  always @(posedge ap_clk) begin
    add_ln160_reg_1586[0] <= 1'b0;
    add_ln160_2_reg_1599[0] <= 1'b0;
    add_ln170_reg_1636[0] <= 1'b0;
    zext_ln52_reg_1641[1:0] <= 2'b00;
    zext_ln52_reg_1641[9] <= 1'b0;
    add_ln52_reg_1646[0] <= 1'b0;
    add_ln21_reg_1680[0] <= 1'b0;
    select_ln40_reg_1685[0] <= 1'b0;
    add_ln23_reg_1690[0] <= 1'b0;
    zext_ln23_2_reg_1703[8:4] <= 5'b00000;
    add_ln112_reg_1754[0] <= 1'b0;
    zext_ln52_3_reg_1775[4] <= 1'b0;
    add_ln73_1_reg_1818[0] <= 1'b0;
    deltas_addr_2_reg_1823[4] <= 1'b0;
    add_ln90_reg_1874[0] <= 1'b0;
    add_ln90_1_reg_1880[0] <= 1'b0;
    select_ln87_reg_1885[0] <= 1'b0;
    add_ln90_3_reg_1915[0] <= 1'b0;
    add_ln90_5_reg_1920[0] <= 1'b0;
  end


endmodule


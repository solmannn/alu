
module reset
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  dec_detl,
  dec_detl_ap_vld,
  detl,
  detl_ap_vld,
  dec_deth,
  dec_deth_ap_vld,
  deth,
  deth_ap_vld,
  rlt2,
  rlt2_ap_vld,
  rlt1,
  rlt1_ap_vld,
  plt2,
  plt2_ap_vld,
  plt1,
  plt1_ap_vld,
  al2,
  al2_ap_vld,
  al1,
  al1_ap_vld,
  nbl,
  nbl_ap_vld,
  rh2,
  rh2_ap_vld,
  rh1,
  rh1_ap_vld,
  ph2,
  ph2_ap_vld,
  ph1,
  ph1_ap_vld,
  ah2,
  ah2_ap_vld,
  ah1,
  ah1_ap_vld,
  nbh,
  nbh_ap_vld,
  dec_rlt2,
  dec_rlt2_ap_vld,
  dec_rlt1,
  dec_rlt1_ap_vld,
  dec_plt2,
  dec_plt2_ap_vld,
  dec_plt1,
  dec_plt1_ap_vld,
  dec_al2,
  dec_al2_ap_vld,
  dec_al1,
  dec_al1_ap_vld,
  dec_nbl,
  dec_nbl_ap_vld,
  dec_rh2,
  dec_rh2_ap_vld,
  dec_rh1,
  dec_rh1_ap_vld,
  dec_ph2,
  dec_ph2_ap_vld,
  dec_ph1,
  dec_ph1_ap_vld,
  dec_ah2,
  dec_ah2_ap_vld,
  dec_ah1,
  dec_ah1_ap_vld,
  dec_nbh,
  dec_nbh_ap_vld,
  delay_dltx_address0,
  delay_dltx_ce0,
  delay_dltx_we0,
  delay_dltx_d0,
  delay_dhx_address0,
  delay_dhx_ce0,
  delay_dhx_we0,
  delay_dhx_d0,
  dec_del_dltx_address0,
  dec_del_dltx_ce0,
  dec_del_dltx_we0,
  dec_del_dltx_d0,
  dec_del_dhx_address0,
  dec_del_dhx_ce0,
  dec_del_dhx_we0,
  dec_del_dhx_d0,
  delay_bpl_address0,
  delay_bpl_ce0,
  delay_bpl_we0,
  delay_bpl_d0,
  delay_bph_address0,
  delay_bph_ce0,
  delay_bph_we0,
  delay_bph_d0,
  dec_del_bpl_address0,
  dec_del_bpl_ce0,
  dec_del_bpl_we0,
  dec_del_bpl_d0,
  dec_del_bph_address0,
  dec_del_bph_ce0,
  dec_del_bph_we0,
  dec_del_bph_d0,
  tqmf_address0,
  tqmf_ce0,
  tqmf_we0,
  tqmf_d0,
  accumc_address0,
  accumc_ce0,
  accumc_we0,
  accumc_d0,
  accumd_address0,
  accumd_ce0,
  accumd_we0,
  accumd_d0,
  working_key
);

  parameter ap_ST_fsm_state1 = 5'd1;
  parameter ap_ST_fsm_state2 = 5'd2;
  parameter ap_ST_fsm_state3 = 5'd4;
  parameter ap_ST_fsm_state4 = 5'd8;
  parameter ap_ST_fsm_state5 = 5'd16;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [14:0] dec_detl;
  output dec_detl_ap_vld;
  output [31:0] detl;
  output detl_ap_vld;
  output [14:0] dec_deth;
  output dec_deth_ap_vld;
  output [14:0] deth;
  output deth_ap_vld;
  output [31:0] rlt2;
  output rlt2_ap_vld;
  output [31:0] rlt1;
  output rlt1_ap_vld;
  output [31:0] plt2;
  output plt2_ap_vld;
  output [31:0] plt1;
  output plt1_ap_vld;
  output [31:0] al2;
  output al2_ap_vld;
  output [31:0] al1;
  output al1_ap_vld;
  output [31:0] nbl;
  output nbl_ap_vld;
  output [31:0] rh2;
  output rh2_ap_vld;
  output [31:0] rh1;
  output rh1_ap_vld;
  output [31:0] ph2;
  output ph2_ap_vld;
  output [31:0] ph1;
  output ph1_ap_vld;
  output [31:0] ah2;
  output ah2_ap_vld;
  output [31:0] ah1;
  output ah1_ap_vld;
  output [31:0] nbh;
  output nbh_ap_vld;
  output [31:0] dec_rlt2;
  output dec_rlt2_ap_vld;
  output [31:0] dec_rlt1;
  output dec_rlt1_ap_vld;
  output [31:0] dec_plt2;
  output dec_plt2_ap_vld;
  output [31:0] dec_plt1;
  output dec_plt1_ap_vld;
  output [31:0] dec_al2;
  output dec_al2_ap_vld;
  output [31:0] dec_al1;
  output dec_al1_ap_vld;
  output [31:0] dec_nbl;
  output dec_nbl_ap_vld;
  output [31:0] dec_rh2;
  output dec_rh2_ap_vld;
  output [31:0] dec_rh1;
  output dec_rh1_ap_vld;
  output [31:0] dec_ph2;
  output dec_ph2_ap_vld;
  output [31:0] dec_ph1;
  output dec_ph1_ap_vld;
  output [31:0] dec_ah2;
  output dec_ah2_ap_vld;
  output [31:0] dec_ah1;
  output dec_ah1_ap_vld;
  output [31:0] dec_nbh;
  output dec_nbh_ap_vld;
  output [2:0] delay_dltx_address0;
  output delay_dltx_ce0;
  output delay_dltx_we0;
  output [31:0] delay_dltx_d0;
  output [2:0] delay_dhx_address0;
  output delay_dhx_ce0;
  output delay_dhx_we0;
  output [31:0] delay_dhx_d0;
  output [2:0] dec_del_dltx_address0;
  output dec_del_dltx_ce0;
  output dec_del_dltx_we0;
  output [31:0] dec_del_dltx_d0;
  output [2:0] dec_del_dhx_address0;
  output dec_del_dhx_ce0;
  output dec_del_dhx_we0;
  output [31:0] dec_del_dhx_d0;
  output [2:0] delay_bpl_address0;
  output delay_bpl_ce0;
  output delay_bpl_we0;
  output [31:0] delay_bpl_d0;
  output [2:0] delay_bph_address0;
  output delay_bph_ce0;
  output delay_bph_we0;
  output [31:0] delay_bph_d0;
  output [2:0] dec_del_bpl_address0;
  output dec_del_bpl_ce0;
  output dec_del_bpl_we0;
  output [31:0] dec_del_bpl_d0;
  output [2:0] dec_del_bph_address0;
  output dec_del_bph_ce0;
  output dec_del_bph_we0;
  output [31:0] dec_del_bph_d0;
  output [4:0] tqmf_address0;
  output tqmf_ce0;
  output tqmf_we0;
  output [6:0] tqmf_d0;
  output [3:0] accumc_address0;
  output accumc_ce0;
  output accumc_we0;
  output [31:0] accumc_d0;
  output [3:0] accumd_address0;
  output accumd_ce0;
  output accumd_we0;
  output [31:0] accumd_d0;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg dec_detl_ap_vld;
  reg detl_ap_vld;
  reg dec_deth_ap_vld;
  reg deth_ap_vld;
  reg rlt2_ap_vld;
  reg rlt1_ap_vld;
  reg plt2_ap_vld;
  reg plt1_ap_vld;
  reg al2_ap_vld;
  reg al1_ap_vld;
  reg nbl_ap_vld;
  reg rh2_ap_vld;
  reg rh1_ap_vld;
  reg ph2_ap_vld;
  reg ph1_ap_vld;
  reg ah2_ap_vld;
  reg ah1_ap_vld;
  reg nbh_ap_vld;
  reg dec_rlt2_ap_vld;
  reg dec_rlt1_ap_vld;
  reg dec_plt2_ap_vld;
  reg dec_plt1_ap_vld;
  reg dec_al2_ap_vld;
  reg dec_al1_ap_vld;
  reg dec_nbl_ap_vld;
  reg dec_rh2_ap_vld;
  reg dec_rh1_ap_vld;
  reg dec_ph2_ap_vld;
  reg dec_ph1_ap_vld;
  reg dec_ah2_ap_vld;
  reg dec_ah1_ap_vld;
  reg dec_nbh_ap_vld;
  reg delay_dltx_ce0;
  reg delay_dltx_we0;
  reg delay_dhx_ce0;
  reg delay_dhx_we0;
  reg dec_del_dltx_ce0;
  reg dec_del_dltx_we0;
  reg dec_del_dhx_ce0;
  reg dec_del_dhx_we0;
  reg delay_bpl_ce0;
  reg delay_bpl_we0;
  reg delay_bph_ce0;
  reg delay_bph_we0;
  reg dec_del_bpl_ce0;
  reg dec_del_bpl_we0;
  reg dec_del_bph_ce0;
  reg dec_del_bph_we0;
  reg tqmf_ce0;
  reg tqmf_we0;
  reg accumc_ce0;
  reg accumc_we0;
  reg accumd_ce0;
  reg accumd_we0;
  reg [4:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  wire [2:0] i_4_fu_520_p2;
  wire ap_CS_fsm_state2;
  wire [2:0] i_5_fu_540_p2;
  wire ap_CS_fsm_state3;
  wire [4:0] i_6_fu_560_p2;
  wire ap_CS_fsm_state4;
  wire [3:0] i_7_fu_577_p2;
  wire ap_CS_fsm_state5;
  reg [2:0] i_reg_278;
  wire [0:0] exitcond3_fu_514_p2;
  reg [2:0] i_1_reg_289;
  wire [0:0] exitcond2_fu_534_p2;
  reg [4:0] i_2_reg_300;
  wire [0:0] exitcond1_fu_554_p2;
  reg [3:0] i_3_reg_311;
  wire [0:0] exitcond_fu_571_p2;
  wire [63:0] tmp_fu_526_p1;
  wire [63:0] tmp_s_fu_546_p1;
  wire [63:0] tmp_11_fu_566_p1;
  wire [63:0] tmp_12_fu_583_p1;
  reg [4:0] ap_NS_fsm;
  input [109:0] working_key;

  initial begin
    #0 ap_CS_fsm = 5'd1;
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state2) & (exitcond3_fu_514_p2 == 1'd1)) begin
      i_1_reg_289 <= 3'd0;
    end else if((exitcond2_fu_534_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3)) begin
      i_1_reg_289 <= i_5_fu_540_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond2_fu_534_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state3)) begin
      i_2_reg_300 <= 5'd0;
    end else if((exitcond1_fu_554_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state4)) begin
      i_2_reg_300 <= i_6_fu_560_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond1_fu_554_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state4)) begin
      i_3_reg_311 <= 4'd0;
    end else if((exitcond_fu_571_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state5)) begin
      i_3_reg_311 <= i_7_fu_577_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state2) & (exitcond3_fu_514_p2 == 1'd0)) begin
      i_reg_278 <= i_4_fu_520_p2;
    end else if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      i_reg_278 <= 3'd0;
    end 
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      accumc_ce0 = 1'b1;
    end else begin
      accumc_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond_fu_571_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state5)) begin
      accumc_we0 = 1'b1;
    end else begin
      accumc_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      accumd_ce0 = 1'b1;
    end else begin
      accumd_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond_fu_571_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state5)) begin
      accumd_we0 = 1'b1;
    end else begin
      accumd_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      ah1_ap_vld = 1'b1;
    end else begin
      ah1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      ah2_ap_vld = 1'b1;
    end else begin
      ah2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      al1_ap_vld = 1'b1;
    end else begin
      al1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      al2_ap_vld = 1'b1;
    end else begin
      al2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond_fu_571_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state5) | (ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond_fu_571_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state5)) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_ah1_ap_vld = 1'b1;
    end else begin
      dec_ah1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_ah2_ap_vld = 1'b1;
    end else begin
      dec_ah2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_al1_ap_vld = 1'b1;
    end else begin
      dec_al1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_al2_ap_vld = 1'b1;
    end else begin
      dec_al2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      dec_del_bph_ce0 = 1'b1;
    end else begin
      dec_del_bph_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond2_fu_534_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3)) begin
      dec_del_bph_we0 = 1'b1;
    end else begin
      dec_del_bph_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      dec_del_bpl_ce0 = 1'b1;
    end else begin
      dec_del_bpl_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond2_fu_534_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3)) begin
      dec_del_bpl_we0 = 1'b1;
    end else begin
      dec_del_bpl_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      dec_del_dhx_ce0 = 1'b1;
    end else begin
      dec_del_dhx_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) & (exitcond3_fu_514_p2 == 1'd0)) begin
      dec_del_dhx_we0 = 1'b1;
    end else begin
      dec_del_dhx_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      dec_del_dltx_ce0 = 1'b1;
    end else begin
      dec_del_dltx_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) & (exitcond3_fu_514_p2 == 1'd0)) begin
      dec_del_dltx_we0 = 1'b1;
    end else begin
      dec_del_dltx_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_deth_ap_vld = 1'b1;
    end else begin
      dec_deth_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_detl_ap_vld = 1'b1;
    end else begin
      dec_detl_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_nbh_ap_vld = 1'b1;
    end else begin
      dec_nbh_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_nbl_ap_vld = 1'b1;
    end else begin
      dec_nbl_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_ph1_ap_vld = 1'b1;
    end else begin
      dec_ph1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_ph2_ap_vld = 1'b1;
    end else begin
      dec_ph2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_plt1_ap_vld = 1'b1;
    end else begin
      dec_plt1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_plt2_ap_vld = 1'b1;
    end else begin
      dec_plt2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_rh1_ap_vld = 1'b1;
    end else begin
      dec_rh1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_rh2_ap_vld = 1'b1;
    end else begin
      dec_rh2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_rlt1_ap_vld = 1'b1;
    end else begin
      dec_rlt1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      dec_rlt2_ap_vld = 1'b1;
    end else begin
      dec_rlt2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      delay_bph_ce0 = 1'b1;
    end else begin
      delay_bph_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond2_fu_534_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3)) begin
      delay_bph_we0 = 1'b1;
    end else begin
      delay_bph_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      delay_bpl_ce0 = 1'b1;
    end else begin
      delay_bpl_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond2_fu_534_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3)) begin
      delay_bpl_we0 = 1'b1;
    end else begin
      delay_bpl_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      delay_dhx_ce0 = 1'b1;
    end else begin
      delay_dhx_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) & (exitcond3_fu_514_p2 == 1'd0)) begin
      delay_dhx_we0 = 1'b1;
    end else begin
      delay_dhx_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      delay_dltx_ce0 = 1'b1;
    end else begin
      delay_dltx_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) & (exitcond3_fu_514_p2 == 1'd0)) begin
      delay_dltx_we0 = 1'b1;
    end else begin
      delay_dltx_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      deth_ap_vld = 1'b1;
    end else begin
      deth_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      detl_ap_vld = 1'b1;
    end else begin
      detl_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      nbh_ap_vld = 1'b1;
    end else begin
      nbh_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      nbl_ap_vld = 1'b1;
    end else begin
      nbl_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      ph1_ap_vld = 1'b1;
    end else begin
      ph1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      ph2_ap_vld = 1'b1;
    end else begin
      ph2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      plt1_ap_vld = 1'b1;
    end else begin
      plt1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      plt2_ap_vld = 1'b1;
    end else begin
      plt2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      rh1_ap_vld = 1'b1;
    end else begin
      rh1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      rh2_ap_vld = 1'b1;
    end else begin
      rh2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      rlt1_ap_vld = 1'b1;
    end else begin
      rlt1_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      rlt2_ap_vld = 1'b1;
    end else begin
      rlt2_ap_vld = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state4) begin
      tqmf_ce0 = 1'b1;
    end else begin
      tqmf_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond1_fu_554_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state4)) begin
      tqmf_we0 = 1'b1;
    end else begin
      tqmf_we0 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if((1'b1 == ap_CS_fsm_state2) & (exitcond3_fu_514_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end
      end
      ap_ST_fsm_state3: begin
        if((exitcond2_fu_534_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state3)) begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end
      end
      ap_ST_fsm_state4: begin
        if((exitcond1_fu_554_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state4)) begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end
      end
      ap_ST_fsm_state5: begin
        if((exitcond_fu_571_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state5)) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign accumc_address0 = tmp_12_fu_583_p1;
  assign accumc_d0 = 32'd0;
  assign accumd_address0 = tmp_12_fu_583_p1;
  assign accumd_d0 = 32'd0;
  assign ah1 = 32'd0;
  assign ah2 = 32'd0;
  assign al1 = 32'd0;
  assign al2 = 32'd0;
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign dec_ah1 = 32'd0;
  assign dec_ah2 = 32'd0;
  assign dec_al1 = 32'd0;
  assign dec_al2 = 32'd0;
  assign dec_del_bph_address0 = tmp_s_fu_546_p1;
  assign dec_del_bph_d0 = 32'd0;
  assign dec_del_bpl_address0 = tmp_s_fu_546_p1;
  assign dec_del_bpl_d0 = 32'd0;
  assign dec_del_dhx_address0 = tmp_fu_526_p1;
  assign dec_del_dhx_d0 = 32'd0;
  assign dec_del_dltx_address0 = tmp_fu_526_p1;
  assign dec_del_dltx_d0 = 32'd0;
  assign dec_deth = 15'd8;
  assign dec_detl = 15'd32;
  assign dec_nbh = 32'd0;
  assign dec_nbl = 32'd0;
  assign dec_ph1 = 32'd0;
  assign dec_ph2 = 32'd0;
  assign dec_plt1 = 32'd0;
  assign dec_plt2 = 32'd0;
  assign dec_rh1 = 32'd0;
  assign dec_rh2 = 32'd0;
  assign dec_rlt1 = 32'd0;
  assign dec_rlt2 = 32'd0;
  assign delay_bph_address0 = tmp_s_fu_546_p1;
  assign delay_bph_d0 = 32'd0;
  assign delay_bpl_address0 = tmp_s_fu_546_p1;
  assign delay_bpl_d0 = 32'd0;
  assign delay_dhx_address0 = tmp_fu_526_p1;
  assign delay_dhx_d0 = 32'd0;
  assign delay_dltx_address0 = tmp_fu_526_p1;
  assign delay_dltx_d0 = 32'd0;
  assign deth = 15'd8;
  assign detl = 32'd32;
  assign exitcond1_fu_554_p2 = (i_2_reg_300 == 5'd24)? 1'b1 : 1'b0;
  assign exitcond2_fu_534_p2 = (i_1_reg_289 == 3'd6)? 1'b1 : 1'b0;
  assign exitcond3_fu_514_p2 = (i_reg_278 == 3'd6)? 1'b1 : 1'b0;
  assign exitcond_fu_571_p2 = (i_3_reg_311 == 4'd11)? 1'b1 : 1'b0;
  assign i_4_fu_520_p2 = i_reg_278 + 3'd1;
  assign i_5_fu_540_p2 = i_1_reg_289 + 3'd1;
  assign i_6_fu_560_p2 = i_2_reg_300 + 5'd1;
  assign i_7_fu_577_p2 = i_3_reg_311 + 4'd1;
  assign nbh = 32'd0;
  assign nbl = 32'd0;
  assign ph1 = 32'd0;
  assign ph2 = 32'd0;
  assign plt1 = 32'd0;
  assign plt2 = 32'd0;
  assign rh1 = 32'd0;
  assign rh2 = 32'd0;
  assign rlt1 = 32'd0;
  assign rlt2 = 32'd0;
  assign tmp_11_fu_566_p1 = i_2_reg_300;
  assign tmp_12_fu_583_p1 = i_3_reg_311;
  assign tmp_fu_526_p1 = i_reg_278;
  assign tmp_s_fu_546_p1 = i_1_reg_289;
  assign tqmf_address0 = tmp_11_fu_566_p1;
  assign tqmf_d0 = 7'd0;

endmodule


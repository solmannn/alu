
module alu
(
  in1,
  in2,
  in3,
  sel,
  out1,
  out2
);

  input [7:0] in1;
  input [7:0] in2;
  input [7:0] in3;
  input sel;
  output [7:0] out1;
  output [7:0] out2;

  alu_0_obf
  i0
  (
    .in1(in1),
    .in2(in2),
    .in3(in3),
    .sel(sel),
    .out1(out1),
    .out2(out2),
    .working_key(255'b110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111)
  );


endmodule



module Gsm_LPC_Analysis_0_obf
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  s_address0,
  s_ce0,
  s_we0,
  s_d0,
  s_q0,
  s_address1,
  s_ce1,
  s_we1,
  s_d1,
  s_q1,
  LARc_address0,
  LARc_ce0,
  LARc_we0,
  LARc_d0,
  LARc_q0,
  LARc_address1,
  LARc_ce1,
  LARc_we1,
  LARc_d1,
  LARc_q1,
  locking_key
);

  parameter ap_ST_fsm_state1 = 60'd1;
  parameter ap_ST_fsm_state2 = 60'd2;
  parameter ap_ST_fsm_state3 = 60'd4;
  parameter ap_ST_fsm_state4 = 60'd8;
  parameter ap_ST_fsm_state5 = 60'd16;
  parameter ap_ST_fsm_state6 = 60'd32;
  parameter ap_ST_fsm_state7 = 60'd64;
  parameter ap_ST_fsm_state8 = 60'd128;
  parameter ap_ST_fsm_state9 = 60'd256;
  parameter ap_ST_fsm_state10 = 60'd512;
  parameter ap_ST_fsm_state11 = 60'd1024;
  parameter ap_ST_fsm_state12 = 60'd2048;
  parameter ap_ST_fsm_state13 = 60'd4096;
  parameter ap_ST_fsm_state14 = 60'd8192;
  parameter ap_ST_fsm_state15 = 60'd16384;
  parameter ap_ST_fsm_state16 = 60'd32768;
  parameter ap_ST_fsm_state17 = 60'd65536;
  parameter ap_ST_fsm_state18 = 60'd131072;
  parameter ap_ST_fsm_state19 = 60'd262144;
  parameter ap_ST_fsm_state20 = 60'd524288;
  parameter ap_ST_fsm_state21 = 60'd1048576;
  parameter ap_ST_fsm_state22 = 60'd2097152;
  parameter ap_ST_fsm_state23 = 60'd4194304;
  parameter ap_ST_fsm_state24 = 60'd8388608;
  parameter ap_ST_fsm_state25 = 60'd16777216;
  parameter ap_ST_fsm_state26 = 60'd33554432;
  parameter ap_ST_fsm_state27 = 60'd67108864;
  parameter ap_ST_fsm_state28 = 60'd134217728;
  parameter ap_ST_fsm_state29 = 60'd268435456;
  parameter ap_ST_fsm_state30 = 60'd536870912;
  parameter ap_ST_fsm_state31 = 60'd1073741824;
  parameter ap_ST_fsm_state32 = 60'd2147483648;
  parameter ap_ST_fsm_state33 = 60'd4294967296;
  parameter ap_ST_fsm_state34 = 60'd8589934592;
  parameter ap_ST_fsm_state35 = 60'd17179869184;
  parameter ap_ST_fsm_state36 = 60'd34359738368;
  parameter ap_ST_fsm_state37 = 60'd68719476736;
  parameter ap_ST_fsm_state38 = 60'd137438953472;
  parameter ap_ST_fsm_state39 = 60'd274877906944;
  parameter ap_ST_fsm_state40 = 60'd549755813888;
  parameter ap_ST_fsm_state41 = 60'd1099511627776;
  parameter ap_ST_fsm_state42 = 60'd2199023255552;
  parameter ap_ST_fsm_state43 = 60'd4398046511104;
  parameter ap_ST_fsm_state44 = 60'd8796093022208;
  parameter ap_ST_fsm_state45 = 60'd17592186044416;
  parameter ap_ST_fsm_state46 = 60'd35184372088832;
  parameter ap_ST_fsm_state47 = 60'd70368744177664;
  parameter ap_ST_fsm_state48 = 60'd140737488355328;
  parameter ap_ST_fsm_state49 = 60'd281474976710656;
  parameter ap_ST_fsm_state50 = 60'd562949953421312;
  parameter ap_ST_fsm_state51 = 60'd1125899906842624;
  parameter ap_ST_fsm_state52 = 60'd2251799813685248;
  parameter ap_ST_fsm_state53 = 60'd4503599627370496;
  parameter ap_ST_fsm_state54 = 60'd9007199254740992;
  parameter ap_ST_fsm_state55 = 60'd18014398509481984;
  parameter ap_ST_fsm_state56 = 60'd36028797018963968;
  parameter ap_ST_fsm_state57 = 60'd72057594037927936;
  parameter ap_ST_fsm_state58 = 60'd144115188075855872;
  parameter ap_ST_fsm_state59 = 60'd288230376151711744;
  parameter ap_ST_fsm_state60 = 60'd576460752303423488;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [7:0] s_address0;
  output s_ce0;
  output s_we0;
  output [15:0] s_d0;
  input [15:0] s_q0;
  output [7:0] s_address1;
  output s_ce1;
  output s_we1;
  output [15:0] s_d1;
  input [15:0] s_q1;
  output [2:0] LARc_address0;
  output LARc_ce0;
  output LARc_we0;
  output [15:0] LARc_d0;
  input [15:0] LARc_q0;
  output [2:0] LARc_address1;
  output LARc_ce1;
  output LARc_we1;
  output [15:0] LARc_d1;
  input [15:0] LARc_q1;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [7:0] s_address0;
  reg s_ce0;
  reg s_we0;
  reg [7:0] s_address1;
  reg s_ce1;
  reg s_we1;
  reg [2:0] LARc_address0;
  reg LARc_ce0;
  reg LARc_we0;
  reg [15:0] LARc_d0;
  reg [2:0] LARc_address1;
  reg LARc_ce1;
  reg LARc_we1;
  reg [15:0] LARc_d1;
  reg [59:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  reg [7:0] bitoff_address0;
  reg bitoff_ce0;
  wire [3:0] bitoff_q0;
  reg [7:0] bitoff_address1;
  reg bitoff_ce1;
  wire [3:0] bitoff_q1;
  reg [7:0] bitoff_address2;
  reg bitoff_ce2;
  wire [3:0] bitoff_q2;
  wire [7:0] bitoff_address3;
  reg bitoff_ce3;
  wire [3:0] bitoff_q3;
  reg [15:0] reg_1099;
  wire ap_CS_fsm_state9;
  wire ap_CS_fsm_state14;
  wire ap_CS_fsm_state21;
  wire [63:0] L_ACF_q0;
  reg [63:0] reg_1104;
  wire ap_CS_fsm_state13;
  wire [63:0] L_ACF_q1;
  wire ap_CS_fsm_state23;
  reg [63:0] reg_1109;
  wire ap_CS_fsm_state15;
  reg [63:0] reg_1114;
  wire ap_CS_fsm_state22;
  wire ap_CS_fsm_state24;
  reg [63:0] reg_1118;
  wire signed [15:0] P_q0;
  reg signed [15:0] reg_1122;
  wire ap_CS_fsm_state43;
  wire ap_CS_fsm_state48;
  wire [7:0] k_fu_1132_p2;
  reg [7:0] k_reg_4621;
  wire ap_CS_fsm_state2;
  wire [0:0] icmp_ln58_fu_1126_p2;
  wire [0:0] icmp_ln118_fu_1151_p2;
  reg [0:0] icmp_ln118_reg_4631;
  wire [0:0] tmp_1_fu_1157_p3;
  reg [0:0] tmp_1_reg_4637;
  wire [0:0] icmp_ln123_fu_1215_p2;
  reg [0:0] icmp_ln123_reg_4642;
  wire [0:0] icmp_ln123_1_fu_1231_p2;
  reg [0:0] icmp_ln123_1_reg_4648;
  wire [0:0] icmp_ln123_2_fu_1286_p2;
  reg [0:0] icmp_ln123_2_reg_4668;
  wire [15:0] select_ln61_fu_1334_p3;
  wire ap_CS_fsm_state3;
  wire signed [15:0] sext_ln67_fu_1479_p1;
  reg signed [15:0] sext_ln67_reg_4678;
  wire ap_CS_fsm_state4;
  wire [0:0] icmp_ln72_fu_1483_p2;
  reg [0:0] icmp_ln72_reg_4683;
  wire [0:0] and_ln72_fu_1495_p2;
  reg [0:0] and_ln72_reg_4687;
  wire [2:0] trunc_ln76_fu_1501_p1;
  reg [2:0] trunc_ln76_reg_4691;
  wire [30:0] zext_ln75_fu_1520_p1;
  reg [30:0] zext_ln75_reg_4696;
  wire ap_CS_fsm_state5;
  wire [7:0] k_1_fu_1530_p2;
  reg [7:0] k_1_reg_4704;
  wire ap_CS_fsm_state6;
  reg [7:0] s_addr_2_reg_4709;
  wire [0:0] icmp_ln75_fu_1524_p2;
  reg [15:0] trunc_ln2_reg_4714;
  wire ap_CS_fsm_state7;
  wire [4:0] k_2_fu_1571_p2;
  wire ap_CS_fsm_state10;
  wire [0:0] tmp_14_fu_1558_p3;
  reg signed [15:0] sl_1_reg_4732;
  wire ap_CS_fsm_state11;
  wire [3:0] L_ACF_addr_1_reg_4748;
  wire ap_CS_fsm_state12;
  reg signed [15:0] sl_2_reg_4754;
  reg signed [15:0] sl_3_reg_4760;
  wire [3:0] L_ACF_addr_2_reg_4776;
  wire [3:0] L_ACF_addr_3_reg_4782;
  reg signed [15:0] sl_4_reg_4788;
  reg signed [15:0] sl_5_reg_4794;
  wire signed [31:0] sext_ln91_fu_1577_p1;
  reg signed [31:0] sext_ln91_reg_4810;
  wire signed [31:0] sext_ln93_1_fu_1584_p1;
  reg signed [31:0] sext_ln93_1_reg_4818;
  wire signed [31:0] mul_ln93_fu_4296_p2;
  reg signed [31:0] mul_ln93_reg_4826;
  wire signed [31:0] mul_ln94_fu_4302_p2;
  reg signed [31:0] mul_ln94_reg_4831;
  wire signed [31:0] sext_ln96_1_fu_1590_p1;
  reg signed [31:0] sext_ln96_1_reg_4836;
  wire signed [31:0] mul_ln98_fu_4308_p2;
  reg signed [31:0] mul_ln98_reg_4844;
  wire signed [16:0] sext_ln100_fu_1593_p1;
  reg signed [16:0] sext_ln100_reg_4849;
  wire signed [31:0] sext_ln100_1_fu_1596_p1;
  reg signed [31:0] sext_ln100_1_reg_4854;
  wire signed [31:0] mul_ln100_fu_4314_p2;
  reg signed [31:0] mul_ln100_reg_4861;
  wire signed [31:0] mul_ln103_fu_4320_p2;
  reg signed [31:0] mul_ln103_reg_4866;
  wire signed [31:0] sext_ln105_1_fu_1599_p1;
  reg signed [31:0] sext_ln105_1_reg_4871;
  wire signed [31:0] mul_ln107_fu_4326_p2;
  reg signed [31:0] mul_ln107_reg_4880;
  wire [3:0] L_ACF_addr_4_reg_4885;
  wire signed [16:0] sext_ln111_fu_1602_p1;
  reg signed [16:0] sext_ln111_reg_4891;
  wire signed [31:0] sext_ln111_1_fu_1605_p1;
  reg signed [31:0] sext_ln111_1_reg_4896;
  wire signed [31:0] mul_ln116_fu_4332_p2;
  reg signed [31:0] mul_ln116_reg_4906;
  wire [3:0] L_ACF_addr_5_reg_4911;
  wire signed [31:0] mul_ln118_fu_4338_p2;
  reg signed [31:0] mul_ln118_reg_4917;
  wire signed [31:0] mul_ln120_fu_4344_p2;
  reg signed [31:0] mul_ln120_reg_4922;
  wire signed [31:0] mul_ln121_fu_4350_p2;
  reg signed [31:0] mul_ln121_reg_4927;
  wire signed [31:0] mul_ln122_fu_4356_p2;
  reg signed [31:0] mul_ln122_reg_4932;
  wire signed [31:0] mul_ln123_fu_4362_p2;
  reg signed [31:0] mul_ln123_reg_4937;
  wire signed [31:0] mul_ln124_fu_4368_p2;
  reg signed [31:0] mul_ln124_reg_4942;
  wire signed [32:0] grp_fu_4374_p3;
  reg signed [32:0] mul_ln127_reg_4947;
  wire signed [32:0] grp_fu_4382_p3;
  reg signed [32:0] mul_ln127_2_reg_4952;
  wire signed [31:0] mul_ln109_fu_4422_p2;
  reg signed [31:0] mul_ln109_reg_4957;
  wire signed [31:0] mul_ln111_fu_4426_p2;
  reg signed [31:0] mul_ln111_reg_4962;
  wire [3:0] L_ACF_addr_6_reg_4967;
  wire signed [32:0] grp_fu_4410_p3;
  reg signed [32:0] add_ln126_2_reg_4973;
  wire [33:0] add_ln126_7_fu_1672_p2;
  reg [33:0] add_ln126_7_reg_4978;
  wire [63:0] add_ln127_fu_1699_p2;
  reg [63:0] add_ln127_reg_4983;
  wire [63:0] add_ln128_fu_1730_p2;
  reg [63:0] add_ln128_reg_4988;
  wire signed [32:0] grp_fu_4416_p3;
  reg signed [32:0] add_ln129_1_reg_4993;
  wire signed [32:0] grp_fu_4437_p3;
  reg signed [32:0] add_ln129_4_reg_4998;
  wire signed [32:0] grp_fu_4442_p3;
  reg signed [32:0] add_ln130_3_reg_5003;
  wire [63:0] add_ln131_fu_1745_p2;
  reg [63:0] add_ln131_reg_5008;
  wire signed [32:0] grp_fu_4497_p3;
  reg signed [32:0] add_ln132_1_reg_5013;
  wire signed [31:0] mul_ln133_fu_4504_p2;
  reg signed [31:0] mul_ln133_reg_5018;
  wire [3:0] L_ACF_addr_7_reg_5023;
  wire [63:0] add_ln126_fu_1775_p2;
  reg [63:0] add_ln126_reg_5029;
  wire ap_CS_fsm_state16;
  wire [63:0] add_ln129_fu_1794_p2;
  reg [63:0] add_ln129_reg_5034;
  wire [63:0] add_ln130_fu_1809_p2;
  reg [63:0] add_ln130_reg_5039;
  wire [63:0] add_ln132_fu_1818_p2;
  reg [63:0] add_ln132_reg_5044;
  wire [63:0] add_ln133_fu_1827_p2;
  reg [63:0] add_ln133_reg_5049;
  wire ap_CS_fsm_state19;
  wire [63:0] sp_0_rec_i_cast_fu_1833_p1;
  reg [63:0] sp_0_rec_i_cast_reg_5060;
  wire ap_CS_fsm_state20;
  reg [7:0] s_addr_10_reg_5065;
  wire [7:0] add_ln138_fu_1854_p2;
  reg [7:0] add_ln138_reg_5073;
  wire [0:0] icmp_ln135_fu_1848_p2;
  wire signed [31:0] sext_ln140_fu_1882_p1;
  reg signed [31:0] sext_ln140_reg_5089;
  wire signed [31:0] mul_ln141_fu_4509_p2;
  reg signed [31:0] mul_ln141_reg_5101;
  wire signed [31:0] mul_ln142_fu_4515_p2;
  reg signed [31:0] mul_ln142_reg_5106;
  wire signed [31:0] mul_ln140_fu_4521_p2;
  reg signed [31:0] mul_ln140_reg_5121;
  wire [63:0] add_ln141_fu_1919_p2;
  reg [63:0] add_ln141_reg_5126;
  wire [63:0] add_ln142_1_fu_1928_p2;
  reg [63:0] add_ln142_1_reg_5131;
  wire signed [31:0] mul_ln143_fu_4525_p2;
  reg signed [31:0] mul_ln143_reg_5136;
  wire signed [31:0] mul_ln144_fu_4530_p2;
  reg signed [31:0] mul_ln144_reg_5141;
  wire [63:0] add_ln140_fu_1971_p2;
  reg [63:0] add_ln140_reg_5156;
  wire [63:0] add_ln143_1_fu_1981_p2;
  reg [63:0] add_ln143_1_reg_5161;
  wire [63:0] add_ln144_1_fu_1990_p2;
  reg [63:0] add_ln144_1_reg_5166;
  wire signed [31:0] mul_ln145_fu_4535_p2;
  reg signed [31:0] mul_ln145_reg_5171;
  wire signed [31:0] mul_ln146_fu_4540_p2;
  reg signed [31:0] mul_ln146_reg_5176;
  wire [63:0] add_ln145_1_fu_2007_p2;
  reg [63:0] add_ln145_1_reg_5191;
  wire ap_CS_fsm_state25;
  wire [63:0] add_ln146_1_fu_2016_p2;
  reg [63:0] add_ln146_1_reg_5196;
  wire signed [31:0] mul_ln147_fu_4545_p2;
  reg signed [31:0] mul_ln147_reg_5201;
  wire signed [31:0] mul_ln148_fu_4550_p2;
  reg signed [31:0] mul_ln148_reg_5206;
  wire [63:0] add_ln147_fu_2033_p2;
  reg [63:0] add_ln147_reg_5211;
  wire ap_CS_fsm_state26;
  wire [63:0] add_ln148_fu_2042_p2;
  reg [63:0] add_ln148_reg_5216;
  reg [3:0] L_ACF_addr_9_reg_5224;
  wire ap_CS_fsm_state29;
  wire [0:0] tmp_15_fu_2052_p3;
  wire [4:0] k_3_fu_2065_p2;
  reg [4:0] k_3_reg_5230;
  reg [7:0] s_addr_19_reg_5235;
  wire ap_CS_fsm_state31;
  wire [7:0] add_ln159_fu_2089_p2;
  reg [7:0] add_ln159_reg_5243;
  wire [0:0] icmp_ln178_fu_2101_p2;
  reg [0:0] icmp_ln178_reg_5248;
  wire ap_CS_fsm_state33;
  wire [0:0] icmp_ln118_1_fu_2107_p2;
  reg [0:0] icmp_ln118_1_reg_5252;
  wire [0:0] sel_tmp57_fu_2321_p2;
  reg [0:0] sel_tmp57_reg_5277;
  wire [0:0] or_ln118_fu_2349_p2;
  reg [0:0] or_ln118_reg_5282;
  wire [0:0] or_ln118_2_fu_2361_p2;
  reg [0:0] or_ln118_2_reg_5287;
  wire signed [31:0] sext_ln187_fu_2439_p1;
  reg signed [31:0] sext_ln187_reg_5292;
  wire ap_CS_fsm_state34;
  wire [3:0] i_fu_2449_p2;
  reg [3:0] i_reg_5300;
  wire ap_CS_fsm_state35;
  wire [63:0] zext_ln187_fu_2455_p1;
  reg [63:0] zext_ln187_reg_5305;
  wire [0:0] icmp_ln186_fu_2443_p2;
  wire [63:0] zext_ln193_fu_2486_p1;
  reg [63:0] zext_ln193_reg_5318;
  wire ap_CS_fsm_state37;
  wire [0:0] icmp_ln192_fu_2480_p2;
  wire [3:0] i_1_fu_2491_p2;
  reg [3:0] i_1_reg_5328;
  wire [3:0] i_2_fu_2503_p2;
  reg [3:0] i_2_reg_5336;
  wire ap_CS_fsm_state39;
  wire [63:0] zext_ln195_fu_2509_p1;
  reg [63:0] zext_ln195_reg_5341;
  wire [0:0] icmp_ln194_fu_2497_p2;
  reg [2:0] LARc_addr_2_reg_5361;
  wire ap_CS_fsm_state42;
  reg signed [15:0] temp_3_reg_5366;
  wire [3:0] add_ln199_fu_2527_p2;
  reg [3:0] add_ln199_reg_5377;
  wire [15:0] zext_ln72_fu_2551_p1;
  wire [0:0] tmp_21_fu_2519_p3;
  wire [0:0] icmp_ln204_fu_2555_p2;
  reg [0:0] icmp_ln204_reg_5387;
  wire signed [63:0] sext_ln138_fu_2561_p1;
  wire signed [63:0] sext_ln139_fu_2565_p1;
  reg signed [63:0] sext_ln139_reg_5396;
  wire signed [16:0] sext_ln139_1_fu_2569_p1;
  reg signed [16:0] sext_ln139_1_reg_5402;
  wire [0:0] icmp_ln147_fu_2573_p2;
  reg [0:0] icmp_ln147_reg_5407;
  wire [4:0] zext_ln206_1_fu_2579_p1;
  reg [4:0] zext_ln206_1_reg_5411;
  wire [3:0] add_ln150_fu_2583_p2;
  wire ap_CS_fsm_state44;
  wire [63:0] L_num_3_fu_2611_p3;
  wire [0:0] icmp_ln150_fu_2589_p2;
  wire [15:0] div_fu_2629_p3;
  wire signed [15:0] select_ln213_fu_2648_p3;
  reg signed [15:0] select_ln213_reg_5434;
  wire [31:0] add_ln207_fu_2683_p2;
  wire [0:0] icmp_ln58_1_fu_2689_p2;
  reg [0:0] icmp_ln58_1_reg_5451;
  wire ap_CS_fsm_state45;
  wire signed [31:0] sext_ln62_2_fu_2703_p1;
  reg signed [31:0] sext_ln62_2_reg_5457;
  wire [15:0] select_ln40_1_fu_2774_p3;
  reg [15:0] select_ln40_1_reg_5463;
  wire [31:0] sub_ln223_fu_2782_p2;
  reg [31:0] sub_ln223_reg_5468;
  wire ap_CS_fsm_state46;
  wire [63:0] zext_ln225_fu_2793_p1;
  reg [63:0] zext_ln225_reg_5476;
  wire ap_CS_fsm_state47;
  wire [0:0] icmp_ln223_fu_2788_p2;
  reg [3:0] K_addr_1_reg_5481;
  wire [31:0] m_fu_2798_p2;
  reg [31:0] m_reg_5486;
  wire [31:0] n_1_fu_2809_p2;
  wire [31:0] add_ln199_2_fu_2815_p2;
  wire signed [15:0] K_q0;
  reg signed [15:0] K_load_reg_5506;
  wire signed [15:0] temp_6_fu_2845_p3;
  reg signed [15:0] temp_6_reg_5512;
  wire signed [15:0] temp_7_fu_2871_p3;
  reg signed [15:0] temp_7_reg_5518;
  wire [3:0] add_ln181_fu_3014_p2;
  wire ap_CS_fsm_state50;
  reg [2:0] LARc_addr_4_reg_5532;
  wire ap_CS_fsm_state51;
  wire [3:0] add_ln253_fu_3031_p2;
  reg [3:0] add_ln253_reg_5541;
  wire [0:0] icmp_ln253_fu_3025_p2;
  wire [15:0] select_ln273_fu_3151_p3;
  reg [15:0] select_ln273_reg_5552;
  wire ap_CS_fsm_state52;
  wire [0:0] icmp_ln40_6_fu_3219_p2;
  reg [0:0] icmp_ln40_6_reg_5557;
  wire ap_CS_fsm_state54;
  reg [6:0] tmp_5_reg_5562;
  wire [0:0] icmp_ln40_7_fu_3301_p2;
  reg [0:0] icmp_ln40_7_reg_5567;
  reg [6:0] tmp_6_reg_5572;
  wire [2:0] LARc_addr_6_reg_5577;
  wire [2:0] LARc_addr_7_reg_5582;
  wire [0:0] icmp_ln40_10_fu_3423_p2;
  reg [0:0] icmp_ln40_10_reg_5587;
  wire ap_CS_fsm_state55;
  reg [6:0] tmp_7_reg_5592;
  wire [0:0] icmp_ln40_8_fu_3495_p2;
  reg [0:0] icmp_ln40_8_reg_5597;
  reg [6:0] tmp_8_reg_5602;
  wire [2:0] LARc_addr_8_reg_5607;
  wire [2:0] LARc_addr_9_reg_5612;
  reg signed [15:0] temp_13_reg_5617;
  wire ap_CS_fsm_state56;
  wire [0:0] icmp_ln40_13_fu_3580_p2;
  reg [0:0] icmp_ln40_13_reg_5623;
  reg [6:0] tmp_s_reg_5628;
  wire [2:0] LARc_addr_10_reg_5633;
  wire [2:0] LARc_addr_11_reg_5638;
  wire [0:0] icmp_ln40_12_fu_3790_p2;
  reg [0:0] icmp_ln40_12_reg_5643;
  wire ap_CS_fsm_state57;
  reg [6:0] tmp_9_reg_5648;
  reg signed [15:0] temp_16_reg_5653;
  reg signed [15:0] temp_17_reg_5659;
  wire [0:0] icmp_ln40_14_fu_3977_p2;
  reg [0:0] icmp_ln40_14_reg_5665;
  wire ap_CS_fsm_state58;
  reg [6:0] tmp_10_reg_5670;
  wire [0:0] icmp_ln40_15_fu_4007_p2;
  reg [0:0] icmp_ln40_15_reg_5675;
  reg [6:0] tmp_11_reg_5680;
  reg [3:0] ACF_address0;
  reg ACF_ce0;
  reg ACF_we0;
  wire [15:0] ACF_d0;
  wire [15:0] ACF_q0;
  reg [3:0] P_address0;
  reg P_ce0;
  reg P_we0;
  reg [15:0] P_d0;
  reg [3:0] K_address0;
  reg K_ce0;
  reg K_we0;
  reg [15:0] K_d0;
  reg [3:0] L_ACF_address0;
  reg L_ACF_ce0;
  reg L_ACF_we0;
  reg [63:0] L_ACF_d0;
  reg [3:0] L_ACF_address1;
  reg L_ACF_ce1;
  reg L_ACF_we1;
  reg [63:0] L_ACF_d1;
  reg [15:0] smax_0_i_reg_839;
  reg [7:0] k_0_i_reg_851;
  reg [7:0] k_1_i_reg_862;
  wire ap_CS_fsm_state8;
  reg signed [4:0] k_2_i_reg_873;
  reg [63:0] empty_57_reg_884;
  wire ap_CS_fsm_state28;
  reg [7:0] sp_0_rec_i_reg_894;
  reg signed [4:0] k_3_i_reg_906;
  wire ap_CS_fsm_state30;
  reg [7:0] p_0_rec_i_reg_917;
  wire ap_CS_fsm_state32;
  reg [3:0] i_1_i_reg_928;
  wire ap_CS_fsm_state36;
  reg [3:0] i_2_i_reg_939;
  wire ap_CS_fsm_state38;
  reg [3:0] i_3_i_reg_950;
  wire ap_CS_fsm_state40;
  reg [31:0] indvars_iv142_reg_961;
  reg [31:0] i_3_reg_973;
  reg [3:0] p_1_rec_i_reg_985;
  reg signed [15:0] temp_24_reg_997;
  reg [63:0] L_num_0_i_i_reg_1006;
  reg [15:0] div_0_i_i_reg_1015;
  reg [3:0] k_0_i_i_reg_1026;
  reg [15:0] ap_phi_mux_p_0_i52_i_phi_fu_1041_p4;
  reg [15:0] p_0_i52_i_reg_1037;
  reg [31:0] p_2_rec_i_reg_1049;
  wire [0:0] icmp_ln206_fu_2677_p2;
  reg [31:0] m_0_i_reg_1060;
  wire ap_CS_fsm_state49;
  reg [3:0] p_0_rec_i1_reg_1071;
  wire [0:0] icmp_ln180_fu_3008_p2;
  reg [3:0] p_0_rec_i16_reg_1082;
  wire [0:0] icmp_ln215_fu_2657_p2;
  wire ap_CS_fsm_state53;
  wire [63:0] zext_ln60_fu_1138_p1;
  wire [63:0] select_ln123_fu_1237_p3;
  wire [63:0] zext_ln123_1_fu_1256_p1;
  wire [63:0] zext_ln123_3_fu_1271_p1;
  wire [63:0] zext_ln76_1_fu_1536_p1;
  wire [63:0] zext_ln89_fu_1566_p1;
  wire [63:0] sum17_cast_fu_1843_p1;
  wire [63:0] zext_ln138_1_fu_1866_p1;
  wire [63:0] zext_ln142_fu_1877_p1;
  wire [63:0] zext_ln143_fu_1900_p1;
  wire [63:0] zext_ln144_fu_1911_p1;
  wire [63:0] zext_ln145_fu_1948_p1;
  wire [63:0] zext_ln146_fu_1959_p1;
  wire [63:0] zext_ln138_fu_1964_p1;
  wire [63:0] zext_ln152_fu_2060_p1;
  wire [63:0] p_0_rec_i_cast_fu_2078_p1;
  wire [63:0] zext_ln123_4_fu_2225_p1;
  wire [63:0] zext_ln123_6_fu_2240_p1;
  wire [63:0] zext_ln123_8_fu_2255_p1;
  wire [63:0] zext_ln123_10_fu_2270_p1;
  wire [63:0] zext_ln206_fu_2514_p1;
  wire [63:0] sum42_cast_fu_2672_p1;
  wire [63:0] zext_ln226_fu_2804_p1;
  wire [63:0] p_0_rec_i1_cast_fu_3003_p1;
  wire [63:0] p_0_rec_i16_cast_fu_3020_p1;
  wire ap_CS_fsm_state17;
  wire ap_CS_fsm_state18;
  wire ap_CS_fsm_state27;
  wire [63:0] shl_ln152_fu_2071_p2;
  wire [15:0] select_ln40_5_fu_2994_p3;
  wire ap_CS_fsm_state41;
  wire [15:0] select_ln40_3_fu_2936_p3;
  wire signed [15:0] sext_ln304_1_fu_3662_p1;
  wire signed [15:0] sext_ln305_1_fu_3727_p1;
  wire signed [15:0] sext_ln306_1_fu_3898_p1;
  wire signed [15:0] sext_ln307_1_fu_3963_p1;
  wire ap_CS_fsm_state59;
  wire signed [15:0] sext_ln309_1_fu_4088_p1;
  wire signed [15:0] sext_ln310_1_fu_4153_p1;
  wire ap_CS_fsm_state60;
  wire signed [15:0] sext_ln311_1_fu_4218_p1;
  wire signed [15:0] sext_ln312_1_fu_4283_p1;
  reg signed [15:0] grp_fu_1093_p0;
  wire [31:0] a_assign_1_fu_1143_p3;
  wire [7:0] trunc_ln116_fu_1181_p1;
  wire [31:0] select_ln116_fu_1165_p3;
  wire [23:0] trunc_ln116_1_fu_1185_p3;
  wire [23:0] select_ln116_1_fu_1173_p3;
  wire [31:0] xor_ln116_fu_1193_p2;
  wire [15:0] tmp_2_fu_1205_p4;
  wire [7:0] tmp_3_fu_1221_p4;
  wire [23:0] xor_ln116_1_fu_1199_p2;
  wire [7:0] trunc_ln123_1_fu_1246_p4;
  wire [7:0] trunc_ln123_2_fu_1261_p4;
  wire [23:0] tmp_4_fu_1276_p4;
  wire [0:0] icmp_ln72_1_fu_1300_p2;
  wire [15:0] sub_ln72_fu_1306_p2;
  wire [0:0] tmp_13_fu_1292_p3;
  wire [15:0] select_ln72_fu_1312_p3;
  wire [15:0] smax_fu_1320_p3;
  wire [0:0] icmp_ln61_fu_1328_p2;
  wire [3:0] add_ln123_fu_1352_p2;
  wire [3:0] add_ln123_1_fu_1362_p2;
  wire [0:0] xor_ln123_fu_1372_p2;
  wire [0:0] xor_ln118_fu_1377_p2;
  wire [0:0] tmp_fu_1382_p2;
  wire [0:0] tmp75_fu_1393_p2;
  wire [0:0] sel_tmp37_fu_1403_p2;
  wire [4:0] zext_ln123_fu_1348_p1;
  wire [4:0] newSel_v_fu_1408_p3;
  wire [4:0] newSel_fu_1416_p2;
  wire [0:0] sel_tmp31_fu_1398_p2;
  wire [0:0] sel_tmp24_fu_1388_p2;
  wire [4:0] zext_ln123_2_fu_1358_p1;
  wire signed [4:0] sext_ln123_fu_1368_p1;
  wire [4:0] newSel112_fu_1432_p3;
  wire [0:0] or_cond_fu_1426_p2;
  wire [5:0] newSel_cast_fu_1422_p1;
  wire signed [5:0] newSel112_cast_fu_1440_p1;
  wire [5:0] newSel114_fu_1444_p3;
  wire [0:0] icmp_ln67_fu_1342_p2;
  wire [0:0] or_ln67_fu_1466_p2;
  wire [5:0] select_ln67_fu_1458_p3;
  wire [5:0] sub_ln70_fu_1452_p2;
  wire signed [5:0] n_fu_1471_p3;
  wire [0:0] icmp_ln72_2_fu_1489_p2;
  wire [2:0] add_ln76_fu_1505_p2;
  wire [14:0] zext_ln76_fu_1510_p1;
  wire [14:0] lshr_ln76_fu_1514_p2;
  wire signed [30:0] grp_fu_4288_p3;
  wire signed [31:0] sext_ln88_fu_1554_p1;
  wire signed [15:0] sext_ln118_1_fu_1612_p0;
  wire signed [15:0] sext_ln126_1_fu_1662_p0;
  wire signed [32:0] grp_fu_4390_p3;
  wire signed [32:0] grp_fu_4397_p3;
  wire signed [33:0] sext_ln126_5_fu_1669_p1;
  wire signed [33:0] sext_ln126_4_fu_1666_p1;
  wire signed [63:0] sext_ln94_fu_1623_p1;
  wire signed [63:0] sext_ln127_1_fu_1684_p1;
  wire [63:0] add_ln127_1_fu_1678_p2;
  wire signed [33:0] grp_fu_4456_p4;
  wire signed [63:0] sext_ln127_6_fu_1696_p1;
  wire [63:0] add_ln127_3_fu_1687_p2;
  wire signed [32:0] grp_fu_4403_p3;
  wire signed [63:0] sext_ln128_1_fu_1705_p1;
  wire signed [32:0] grp_fu_4430_p3;
  wire signed [32:0] grp_fu_4465_p3;
  wire signed [33:0] sext_ln128_3_fu_1717_p1;
  wire signed [33:0] sext_ln128_2_fu_1714_p1;
  wire [33:0] add_ln128_5_fu_1720_p2;
  wire signed [63:0] sext_ln128_4_fu_1726_p1;
  wire [63:0] add_ln128_2_fu_1708_p2;
  wire signed [63:0] sext_ln116_fu_1641_p1;
  wire signed [32:0] grp_fu_4489_p3;
  wire signed [63:0] sext_ln131_1_fu_1742_p1;
  wire [63:0] add_ln131_1_fu_1736_p2;
  wire signed [63:0] sext_ln111_2_fu_1754_p1;
  wire signed [63:0] sext_ln126_3_fu_1763_p1;
  wire [63:0] add_ln126_1_fu_1757_p2;
  wire signed [63:0] sext_ln126_6_fu_1772_p1;
  wire [63:0] add_ln126_3_fu_1766_p2;
  wire signed [63:0] sext_ln129_1_fu_1782_p1;
  wire signed [63:0] sext_ln129_2_fu_1791_p1;
  wire [63:0] add_ln129_2_fu_1785_p2;
  wire signed [63:0] sext_ln109_fu_1751_p1;
  wire signed [63:0] sext_ln130_1_fu_1806_p1;
  wire [63:0] add_ln130_1_fu_1800_p2;
  wire signed [63:0] sext_ln132_1_fu_1815_p1;
  wire signed [63:0] sext_ln133_fu_1824_p1;
  wire [7:0] sum17_fu_1837_p2;
  wire [7:0] add_ln138_1_fu_1860_p2;
  wire [7:0] add_ln142_fu_1871_p2;
  wire [7:0] add_ln143_fu_1894_p2;
  wire [7:0] add_ln144_fu_1905_p2;
  wire signed [63:0] sext_ln141_1_fu_1916_p1;
  wire signed [63:0] sext_ln142_1_fu_1925_p1;
  wire [7:0] add_ln145_fu_1942_p2;
  wire [7:0] add_ln146_fu_1953_p2;
  wire signed [63:0] sext_ln140_1_fu_1968_p1;
  wire signed [63:0] sext_ln143_1_fu_1978_p1;
  wire signed [63:0] sext_ln144_1_fu_1987_p1;
  wire signed [63:0] sext_ln145_1_fu_2004_p1;
  wire signed [63:0] sext_ln146_1_fu_2013_p1;
  wire signed [63:0] sext_ln147_1_fu_2030_p1;
  wire signed [63:0] sext_ln148_1_fu_2039_p1;
  wire signed [31:0] sext_ln151_fu_2048_p1;
  wire [0:0] tmp_16_fu_2113_p3;
  wire [7:0] trunc_ln116_5_fu_2165_p1;
  wire [7:0] select_ln116_5_fu_2157_p3;
  wire [15:0] trunc_ln116_4_fu_2153_p1;
  wire [15:0] select_ln116_4_fu_2145_p3;
  wire [31:0] trunc_ln116_2_fu_2129_p1;
  wire [31:0] select_ln116_2_fu_2121_p3;
  wire [23:0] trunc_ln116_3_fu_2141_p1;
  wire [23:0] select_ln116_3_fu_2133_p3;
  wire [31:0] xor_ln95_2_fu_2181_p2;
  wire [15:0] tmp_17_fu_2193_p4;
  wire [7:0] tmp_18_fu_2209_p4;
  wire [7:0] xor_ln95_fu_2169_p2;
  wire [15:0] xor_ln95_1_fu_2175_p2;
  wire [7:0] trunc_ln123_3_fu_2230_p4;
  wire [23:0] xor_ln95_3_fu_2187_p2;
  wire [7:0] trunc_ln123_4_fu_2245_p4;
  wire [7:0] trunc_ln123_5_fu_2260_p4;
  wire [0:0] icmp_ln123_3_fu_2203_p2;
  wire [0:0] xor_ln123_1_fu_2275_p2;
  wire [0:0] xor_ln118_1_fu_2281_p2;
  wire [0:0] tmp110_fu_2287_p2;
  wire [0:0] icmp_ln123_4_fu_2219_p2;
  wire [7:0] tmp_19_fu_2299_p4;
  wire [0:0] icmp_ln123_5_fu_2309_p2;
  wire [0:0] tmp111_fu_2315_p2;
  wire [23:0] tmp_20_fu_2327_p4;
  wire [0:0] icmp_ln123_6_fu_2337_p2;
  wire [0:0] sel_tmp63_fu_2343_p2;
  wire [0:0] sel_tmp50_fu_2293_p2;
  wire [0:0] or_ln118_1_fu_2355_p2;
  wire [4:0] zext_ln123_5_fu_2367_p1;
  wire [4:0] zext_ln123_7_fu_2377_p1;
  wire [3:0] add_ln123_4_fu_2387_p2;
  wire [3:0] add_ln123_5_fu_2397_p2;
  wire [4:0] add_ln123_2_fu_2371_p2;
  wire [4:0] add_ln123_3_fu_2381_p2;
  wire [4:0] zext_ln123_9_fu_2393_p1;
  wire [4:0] select_ln118_fu_2407_p3;
  wire [4:0] select_ln118_1_fu_2414_p3;
  wire [4:0] select_ln118_2_fu_2421_p3;
  wire [5:0] zext_ln118_fu_2428_p1;
  wire signed [5:0] sext_ln123_2_fu_2403_p1;
  wire [5:0] temp_2_fu_2432_p3;
  wire [31:0] trunc_ln187_fu_2460_p1;
  wire [31:0] shl_ln187_fu_2464_p2;
  wire signed [15:0] tmp_21_fu_2519_p1;
  wire signed [15:0] trunc_ln72_fu_2533_p0;
  wire [14:0] trunc_ln72_fu_2533_p1;
  wire [0:0] grp_fu_1093_p2;
  wire [14:0] sub_ln72_1_fu_2537_p2;
  wire [14:0] select_ln72_1_fu_2543_p3;
  wire signed [15:0] icmp_ln204_fu_2555_p0;
  wire signed [15:0] sext_ln139_fu_2565_p0;
  wire signed [15:0] sext_ln139_1_fu_2569_p0;
  wire [63:0] L_num_1_fu_2595_p2;
  wire [0:0] icmp_ln155_fu_2601_p2;
  wire [63:0] L_num_2_fu_2606_p2;
  wire [14:0] trunc_ln155_fu_2625_p1;
  wire [0:0] xor_ln155_fu_2619_p2;
  wire [0:0] icmp_ln213_fu_2637_p2;
  wire [15:0] sub_ln214_fu_2642_p2;
  wire [4:0] empty_65_fu_2663_p1;
  wire [4:0] sum42_fu_2667_p2;
  wire signed [31:0] grp_fu_4555_p3;
  wire [0:0] and_ln58_fu_2694_p2;
  wire [15:0] trunc_ln64_1_fu_2706_p4;
  wire signed [15:0] temp_5_fu_2715_p3;
  wire signed [16:0] sext_ln39_fu_2723_p1;
  wire [16:0] sum_fu_2727_p2;
  wire [1:0] tmp_22_fu_2738_p4;
  wire [0:0] icmp_ln40_fu_2732_p2;
  wire [0:0] icmp_ln40_1_fu_2748_p2;
  wire [0:0] or_ln40_fu_2768_p2;
  wire [15:0] select_ln40_fu_2760_p3;
  wire [15:0] add_ln40_1_fu_2754_p2;
  wire signed [15:0] icmp_ln58_3_fu_2821_p0;
  wire [0:0] icmp_ln58_3_fu_2821_p2;
  wire signed [31:0] grp_fu_4564_p3;
  wire [0:0] and_ln58_1_fu_2827_p2;
  wire [15:0] trunc_ln64_2_fu_2836_p4;
  wire signed [31:0] grp_fu_4572_p3;
  wire [0:0] and_ln58_2_fu_2857_p2;
  wire [15:0] trunc_ln64_3_fu_2862_p4;
  wire signed [16:0] sext_ln39_2_fu_2882_p1;
  wire signed [16:0] sext_ln39_3_fu_2886_p1;
  wire [16:0] sum_1_fu_2889_p2;
  wire [1:0] tmp_23_fu_2901_p4;
  wire [0:0] icmp_ln40_2_fu_2895_p2;
  wire [0:0] icmp_ln40_3_fu_2911_p2;
  wire [0:0] or_ln40_1_fu_2930_p2;
  wire [15:0] select_ln40_2_fu_2922_p3;
  wire [15:0] add_ln40_6_fu_2917_p2;
  wire signed [16:0] sext_ln62_3_fu_2879_p1;
  wire signed [16:0] sext_ln39_4_fu_2945_p1;
  wire [16:0] sum_2_fu_2948_p2;
  wire [1:0] tmp_24_fu_2960_p4;
  wire [0:0] icmp_ln40_4_fu_2954_p2;
  wire [0:0] icmp_ln40_5_fu_2970_p2;
  wire [0:0] or_ln40_2_fu_2988_p2;
  wire [15:0] select_ln40_4_fu_2980_p3;
  wire [15:0] add_ln40_10_fu_2976_p2;
  wire [0:0] icmp_ln72_4_fu_3045_p2;
  wire [15:0] sub_ln72_2_fu_3051_p2;
  wire [0:0] tmp_39_fu_3037_p3;
  wire [15:0] select_ln72_2_fu_3057_p3;
  wire [15:0] temp_fu_3065_p3;
  wire [14:0] trunc_ln5_fu_3079_p4;
  wire [15:0] shl_ln270_fu_3105_p2;
  wire [0:0] icmp_ln259_fu_3073_p2;
  wire signed [15:0] temp_19_fu_3089_p1;
  wire [15:0] temp_21_fu_3111_p2;
  wire [0:0] icmp_ln263_fu_3093_p2;
  wire [0:0] xor_ln259_fu_3125_p2;
  wire [0:0] and_ln263_fu_3131_p2;
  wire [15:0] temp_20_fu_3099_p2;
  wire [15:0] temp_22_fu_3117_p3;
  wire [15:0] temp_23_fu_3137_p3;
  wire [15:0] sub_ln273_fu_3145_p2;
  wire [29:0] shl_ln1_fu_3159_p3;
  wire [27:0] shl_ln50_1_fu_3171_p3;
  wire signed [30:0] sext_ln50_1_fu_3179_p1;
  wire signed [30:0] sext_ln50_fu_3167_p1;
  wire [30:0] add_ln50_fu_3183_p2;
  wire signed [15:0] temp_8_fu_3189_p4;
  wire signed [16:0] sext_ln39_5_fu_3199_p1;
  wire [16:0] sum_3_fu_3203_p2;
  wire [1:0] tmp_25_fu_3209_p4;
  wire [15:0] add_ln40_fu_3225_p2;
  wire [29:0] shl_ln50_2_fu_3241_p3;
  wire [27:0] shl_ln50_3_fu_3253_p3;
  wire signed [30:0] sext_ln50_3_fu_3261_p1;
  wire signed [30:0] sext_ln50_2_fu_3249_p1;
  wire [30:0] add_ln50_1_fu_3265_p2;
  wire signed [15:0] temp_9_fu_3271_p4;
  wire signed [16:0] sext_ln39_6_fu_3281_p1;
  wire [16:0] sum_4_fu_3285_p2;
  wire [1:0] tmp_27_fu_3291_p4;
  wire [15:0] add_ln40_2_fu_3307_p2;
  wire [29:0] shl_ln50_4_fu_3323_p3;
  wire [27:0] shl_ln50_5_fu_3335_p3;
  wire signed [30:0] sext_ln50_5_fu_3343_p1;
  wire signed [30:0] sext_ln50_4_fu_3331_p1;
  wire [30:0] add_ln50_2_fu_3347_p2;
  wire signed [15:0] temp_10_fu_3353_p4;
  wire signed [16:0] sext_ln39_7_fu_3363_p1;
  wire [16:0] sum_5_fu_3367_p2;
  wire [1:0] tmp_29_fu_3373_p4;
  wire [0:0] icmp_ln40_9_fu_3383_p2;
  wire [15:0] add_ln40_3_fu_3389_p2;
  wire signed [15:0] temp_11_fu_3395_p3;
  wire signed [16:0] sext_ln39_8_fu_3403_p1;
  wire [16:0] sum_6_fu_3407_p2;
  wire [1:0] tmp_30_fu_3413_p4;
  wire [15:0] add_ln40_4_fu_3429_p2;
  wire [29:0] shl_ln50_6_fu_3445_p3;
  wire [27:0] shl_ln50_7_fu_3457_p3;
  wire signed [30:0] sext_ln50_7_fu_3465_p1;
  wire signed [30:0] sext_ln50_6_fu_3453_p1;
  wire [30:0] add_ln50_3_fu_3469_p2;
  wire signed [15:0] temp_12_fu_3475_p4;
  wire signed [16:0] sext_ln39_9_fu_3485_p1;
  wire [16:0] sum_7_fu_3489_p2;
  wire [15:0] add_ln40_5_fu_3501_p2;
  wire signed [30:0] mul_ln50_fu_4580_p2;
  wire [29:0] shl_ln50_8_fu_3530_p3;
  wire [25:0] shl_ln50_9_fu_3542_p3;
  wire signed [30:0] sext_ln50_9_fu_3538_p1;
  wire signed [30:0] sext_ln50_10_fu_3550_p1;
  wire [30:0] sub_ln50_fu_3554_p2;
  wire signed [15:0] temp_15_fu_3560_p4;
  wire signed [16:0] sext_ln39_12_fu_3570_p1;
  wire [16:0] sum_10_fu_3574_p2;
  wire [15:0] add_ln40_9_fu_3586_p2;
  wire signed [6:0] select_ln40_6_fu_3602_p3;
  wire [1:0] tmp_26_fu_3612_p4;
  wire signed [7:0] sext_ln304_fu_3608_p1;
  wire [0:0] icmp_ln304_fu_3622_p2;
  wire [0:0] icmp_ln304_1_fu_3628_p2;
  wire [0:0] or_ln304_fu_3648_p2;
  wire [7:0] select_ln304_fu_3640_p3;
  wire [7:0] add_ln304_fu_3634_p2;
  wire [7:0] select_ln304_1_fu_3654_p3;
  wire signed [6:0] select_ln40_7_fu_3667_p3;
  wire [1:0] tmp_28_fu_3677_p4;
  wire signed [7:0] sext_ln305_fu_3673_p1;
  wire [0:0] icmp_ln305_fu_3687_p2;
  wire [0:0] icmp_ln305_1_fu_3693_p2;
  wire [0:0] or_ln305_fu_3713_p2;
  wire [7:0] select_ln305_fu_3705_p3;
  wire [7:0] add_ln305_fu_3699_p2;
  wire [7:0] select_ln305_1_fu_3719_p3;
  wire signed [16:0] sext_ln39_10_fu_3732_p1;
  wire [16:0] sum_8_fu_3735_p2;
  wire [1:0] tmp_33_fu_3741_p4;
  wire [0:0] icmp_ln40_11_fu_3751_p2;
  wire [15:0] add_ln40_7_fu_3757_p2;
  wire signed [15:0] temp_14_fu_3762_p3;
  wire signed [16:0] sext_ln39_11_fu_3770_p1;
  wire [16:0] sum_9_fu_3774_p2;
  wire [1:0] tmp_34_fu_3780_p4;
  wire [15:0] add_ln40_8_fu_3796_p2;
  wire signed [30:0] mul_ln50_1_fu_4587_p2;
  wire signed [30:0] mul_ln50_2_fu_4594_p2;
  wire signed [6:0] select_ln40_9_fu_3838_p3;
  wire [2:0] tmp_31_fu_3848_p4;
  wire signed [7:0] sext_ln306_fu_3844_p1;
  wire [0:0] icmp_ln306_fu_3858_p2;
  wire [0:0] icmp_ln306_1_fu_3864_p2;
  wire [0:0] or_ln306_fu_3884_p2;
  wire [7:0] select_ln306_fu_3876_p3;
  wire [7:0] add_ln306_fu_3870_p2;
  wire [7:0] select_ln306_1_fu_3890_p3;
  wire signed [6:0] select_ln40_10_fu_3903_p3;
  wire [2:0] tmp_32_fu_3913_p4;
  wire signed [7:0] sext_ln307_fu_3909_p1;
  wire [0:0] icmp_ln307_fu_3923_p2;
  wire [0:0] icmp_ln307_1_fu_3929_p2;
  wire [0:0] or_ln307_fu_3949_p2;
  wire [7:0] select_ln307_fu_3941_p3;
  wire [7:0] add_ln307_fu_3935_p2;
  wire [7:0] select_ln307_1_fu_3955_p3;
  wire signed [16:0] sext_ln39_13_fu_3968_p1;
  wire [16:0] sum_11_fu_3971_p2;
  wire [15:0] add_ln40_11_fu_3983_p2;
  wire signed [16:0] sext_ln39_14_fu_3998_p1;
  wire [16:0] sum_12_fu_4001_p2;
  wire [15:0] add_ln40_12_fu_4013_p2;
  wire signed [6:0] select_ln40_12_fu_4028_p3;
  wire [3:0] tmp_35_fu_4038_p4;
  wire signed [7:0] sext_ln309_fu_4034_p1;
  wire [0:0] icmp_ln309_fu_4048_p2;
  wire [0:0] icmp_ln309_1_fu_4054_p2;
  wire [0:0] or_ln309_fu_4074_p2;
  wire [7:0] select_ln309_fu_4066_p3;
  wire [7:0] add_ln309_fu_4060_p2;
  wire [7:0] select_ln309_1_fu_4080_p3;
  wire signed [6:0] select_ln40_13_fu_4093_p3;
  wire [3:0] tmp_36_fu_4103_p4;
  wire signed [7:0] sext_ln310_fu_4099_p1;
  wire [0:0] icmp_ln310_fu_4113_p2;
  wire [0:0] icmp_ln310_1_fu_4119_p2;
  wire [0:0] or_ln310_fu_4139_p2;
  wire [7:0] select_ln310_fu_4131_p3;
  wire [7:0] add_ln310_fu_4125_p2;
  wire [7:0] select_ln310_1_fu_4145_p3;
  wire signed [6:0] select_ln40_14_fu_4158_p3;
  wire [4:0] tmp_37_fu_4168_p4;
  wire signed [7:0] sext_ln311_fu_4164_p1;
  wire [0:0] icmp_ln311_fu_4178_p2;
  wire [0:0] icmp_ln311_1_fu_4184_p2;
  wire [0:0] or_ln311_fu_4204_p2;
  wire [7:0] select_ln311_fu_4196_p3;
  wire [7:0] add_ln311_fu_4190_p2;
  wire [7:0] select_ln311_1_fu_4210_p3;
  wire signed [6:0] select_ln40_15_fu_4223_p3;
  wire [4:0] tmp_38_fu_4233_p4;
  wire signed [7:0] sext_ln312_fu_4229_p1;
  wire [0:0] icmp_ln312_fu_4243_p2;
  wire [0:0] icmp_ln312_1_fu_4249_p2;
  wire [0:0] or_ln312_fu_4269_p2;
  wire [7:0] select_ln312_fu_4261_p3;
  wire [7:0] add_ln312_fu_4255_p2;
  wire [7:0] select_ln312_1_fu_4275_p3;
  wire [14:0] grp_fu_4288_p0;
  wire [15:0] grp_fu_4288_p2;
  wire signed [15:0] mul_ln93_fu_4296_p0;
  wire signed [15:0] mul_ln93_fu_4296_p1;
  wire signed [15:0] mul_ln94_fu_4302_p0;
  wire signed [15:0] mul_ln94_fu_4302_p1;
  wire signed [15:0] mul_ln98_fu_4308_p0;
  wire signed [15:0] mul_ln98_fu_4308_p1;
  wire signed [15:0] mul_ln100_fu_4314_p0;
  wire signed [15:0] mul_ln100_fu_4314_p1;
  wire signed [15:0] mul_ln103_fu_4320_p0;
  wire signed [15:0] mul_ln103_fu_4320_p1;
  wire signed [15:0] mul_ln107_fu_4326_p0;
  wire signed [15:0] mul_ln107_fu_4326_p1;
  wire signed [15:0] mul_ln116_fu_4332_p1;
  wire signed [15:0] mul_ln118_fu_4338_p0;
  wire signed [31:0] sext_ln118_1_fu_1612_p1;
  wire signed [15:0] mul_ln118_fu_4338_p1;
  wire signed [15:0] mul_ln120_fu_4344_p0;
  wire signed [15:0] mul_ln120_fu_4344_p1;
  wire signed [15:0] mul_ln121_fu_4350_p0;
  wire signed [15:0] mul_ln121_fu_4350_p1;
  wire signed [15:0] mul_ln122_fu_4356_p0;
  wire signed [15:0] mul_ln122_fu_4356_p1;
  wire signed [15:0] mul_ln123_fu_4362_p0;
  wire signed [15:0] mul_ln123_fu_4362_p1;
  wire signed [15:0] mul_ln124_fu_4368_p0;
  wire signed [15:0] mul_ln124_fu_4368_p1;
  wire signed [15:0] grp_fu_4390_p0;
  wire signed [15:0] grp_fu_4390_p1;
  wire signed [15:0] grp_fu_4397_p0;
  wire signed [15:0] grp_fu_4397_p1;
  wire signed [32:0] grp_fu_4447_p3;
  wire signed [15:0] grp_fu_4403_p0;
  wire signed [15:0] grp_fu_4403_p1;
  wire signed [15:0] grp_fu_4410_p0;
  wire signed [15:0] grp_fu_4410_p1;
  wire signed [15:0] grp_fu_4416_p0;
  wire signed [15:0] grp_fu_4416_p1;
  wire signed [15:0] mul_ln109_fu_4422_p0;
  wire signed [15:0] mul_ln109_fu_4422_p1;
  wire signed [15:0] mul_ln111_fu_4426_p0;
  wire signed [15:0] mul_ln111_fu_4426_p1;
  wire signed [15:0] grp_fu_4430_p0;
  wire signed [15:0] grp_fu_4430_p1;
  wire signed [15:0] grp_fu_4437_p0;
  wire signed [15:0] grp_fu_4437_p1;
  wire signed [32:0] grp_fu_4473_p3;
  wire signed [15:0] grp_fu_4442_p0;
  wire signed [15:0] grp_fu_4442_p1;
  wire signed [32:0] grp_fu_4481_p3;
  wire signed [15:0] grp_fu_4447_p0;
  wire signed [31:0] sext_ln126_1_fu_1662_p1;
  wire signed [15:0] grp_fu_4447_p1;
  wire signed [15:0] grp_fu_4456_p0;
  wire signed [15:0] grp_fu_4456_p1;
  wire signed [15:0] grp_fu_4465_p0;
  wire signed [15:0] grp_fu_4465_p1;
  wire signed [15:0] grp_fu_4473_p0;
  wire signed [15:0] grp_fu_4473_p1;
  wire signed [15:0] grp_fu_4481_p0;
  wire signed [15:0] grp_fu_4481_p1;
  wire signed [15:0] grp_fu_4489_p0;
  wire signed [15:0] grp_fu_4489_p1;
  wire signed [15:0] grp_fu_4497_p0;
  wire signed [15:0] grp_fu_4497_p1;
  wire signed [15:0] mul_ln133_fu_4504_p0;
  wire signed [15:0] mul_ln133_fu_4504_p1;
  wire signed [15:0] mul_ln141_fu_4509_p1;
  wire signed [15:0] mul_ln142_fu_4515_p1;
  wire signed [15:0] mul_ln140_fu_4521_p0;
  wire signed [15:0] mul_ln140_fu_4521_p1;
  wire signed [15:0] mul_ln143_fu_4525_p1;
  wire signed [15:0] mul_ln144_fu_4530_p1;
  wire signed [15:0] mul_ln145_fu_4535_p1;
  wire signed [15:0] mul_ln146_fu_4540_p1;
  wire signed [15:0] mul_ln147_fu_4545_p1;
  wire signed [15:0] mul_ln148_fu_4550_p1;
  wire [15:0] grp_fu_4555_p2;
  wire signed [15:0] grp_fu_4564_p1;
  wire [15:0] grp_fu_4564_p2;
  wire signed [15:0] grp_fu_4572_p0;
  wire [15:0] grp_fu_4572_p2;
  wire [14:0] mul_ln50_fu_4580_p1;
  wire [14:0] mul_ln50_1_fu_4587_p1;
  wire [14:0] mul_ln50_2_fu_4594_p1;
  wire [0:0] icmp_ln158_fu_2083_p2;
  reg [59:0] ap_NS_fsm;
  wire Const_16;
  wire Const_17;
  wire Const_18;
  wire Const_19;
  wire Const_20;
  wire Const_21;
  wire Const_22;
  wire Const_23;
  wire Const_24;
  wire Const_25;
  wire Const_26;
  wire [15:0] Const_27;
  wire Const_28;
  wire Const_29;
  wire Const_30;
  wire Const_31;
  wire Const_32;
  wire Const_33;
  wire Const_34;
  wire Const_35;
  wire Const_36;
  wire [3:0] Const_37;
  wire Const_38;
  wire Const_39;
  wire [3:0] Const_40;
  wire Const_41;
  wire Const_42;
  wire Const_43;
  wire [3:0] Const_44;
  wire Const_45;
  wire Const_46;
  wire Const_47;
  wire [31:0] Const_48;
  wire Const_49;
  wire Const_50;
  wire Const_51;
  wire Const_52;
  wire [31:0] Const_53;
  wire Const_54;
  wire Const_55;
  wire Const_56;
  wire Const_57;
  wire Const_58;
  wire [3:0] Const_59;
  wire Const_60;
  wire Const_61;
  wire Const_62;
  wire Const_63;
  wire Const_64;
  wire Const_65;
  wire Const_66;
  wire Const_67;
  wire [7:0] Const_68;
  wire Const_69;
  wire [7:0] Const_70;
  wire Const_71;
  wire Const_72;
  wire Const_73;
  wire Const_74;
  wire [4:0] Const_75;
  wire Const_76;
  wire Const_77;
  wire [4:0] Const_78;
  wire Const_79;
  wire Const_80;
  wire Const_81;
  wire [31:0] Const_82;
  wire Const_83;
  wire Const_84;
  wire Const_85;
  wire Const_86;
  wire Const_87;
  wire Const_88;
  wire Const_89;
  wire Const_90;
  wire [15:0] Const_91;
  wire Const_92;
  wire Const_93;
  wire Const_94;
  wire Const_95;
  wire Const_96;
  wire Const_97;
  wire Const_98;
  wire Const_99;
  wire Const_100;
  wire Const_101;
  wire Const_102;
  wire [3:0] Const_103;
  wire Const_104;
  wire Const_105;
  wire [3:0] Const_106;
  wire Const_107;
  wire Const_108;
  wire Const_109;
  wire Const_110;
  wire Const_111;
  wire [7:0] Const_112;
  wire Const_113;
  wire Const_114;
  wire Const_115;
  wire [3:0] Const_116;
  wire Const_117;
  wire Const_118;
  wire Const_119;
  wire Const_120;
  wire [31:0] Const_121;
  wire Const_122;
  wire Const_123;
  wire Const_124;
  wire Const_125;
  wire Const_126;
  wire Const_127;
  wire Const_128;
  wire Const_129;
  wire Const_130;
  wire Const_131;
  wire Const_132;
  wire Const_133;
  wire Const_134;
  wire Const_135;
  wire Const_136;
  wire Const_137;
  wire Const_138;
  wire [15:0] Const_139;
  wire Const_140;
  wire Const_141;
  wire [7:0] Const_142;
  wire Const_143;
  wire Const_144;
  wire Const_145;
  wire Const_146;
  wire Const_147;
  wire Const_148;
  wire Const_149;
  wire Const_150;
  wire Const_151;
  wire Const_152;
  wire Const_153;
  wire Const_154;
  wire Const_155;
  wire Const_156;
  wire Const_157;
  wire Const_158;
  wire Const_159;
  wire Const_160;
  wire Const_161;
  wire Const_162;
  wire Const_163;
  wire Const_164;
  wire Const_165;
  wire Const_166;
  wire Const_167;
  wire Const_168;
  wire Const_169;
  wire Const_170;
  wire Const_171;
  wire Const_172;
  wire Const_173;
  wire Const_174;
  wire Const_175;
  wire Const_176;
  wire Const_177;
  wire Const_178;
  wire Const_179;
  wire Const_180;
  wire Const_181;
  wire Const_182;
  wire Const_183;
  wire Const_184;
  wire Const_185;
  wire Const_186;
  wire Const_187;
  wire Const_188;
  wire Const_189;
  wire Const_190;
  wire Const_191;
  wire Const_192;
  wire Const_193;
  wire Const_194;
  wire Const_195;
  wire Const_196;
  wire Const_197;
  wire Const_198;
  wire Const_199;
  wire Const_200;
  wire Const_201;
  wire Const_202;
  wire Const_203;
  wire Const_204;
  wire Const_205;
  wire Const_206;
  wire Const_207;
  wire Const_208;
  wire Const_209;
  wire Const_210;
  wire Const_211;
  wire Const_212;
  wire Const_213;
  wire Const_214;
  wire Const_215;
  wire Const_216;
  wire Const_217;
  wire Const_218;
  wire Const_219;
  wire Const_220;
  wire Const_221;
  wire Const_222;
  wire Const_223;
  wire Const_224;
  wire Const_225;
  wire Const_226;
  wire Const_227;
  wire Const_228;
  wire Const_229;
  wire Const_230;
  wire Const_231;
  wire Const_232;
  wire Const_233;
  wire Const_234;
  wire Const_235;
  wire Const_236;
  wire Const_237;
  wire Const_238;
  wire Const_239;
  wire Const_240;
  wire Const_241;
  wire Const_242;
  wire Const_243;
  wire Const_244;
  wire Const_245;
  wire [2:0] Const_246;
  wire Const_247;
  wire [2:0] Const_248;
  wire Const_249;
  wire [2:0] Const_250;
  wire Const_251;
  wire [2:0] Const_252;
  wire Const_253;
  wire Const_254;
  wire [2:0] Const_255;
  wire Const_256;
  wire Const_257;
  wire Const_258;
  wire Const_259;
  wire Const_260;
  wire Const_261;
  wire Const_262;
  wire Const_263;
  wire Const_264;
  wire Const_265;
  wire Const_266;
  wire Const_267;
  wire Const_268;
  wire Const_269;
  wire Const_270;
  wire Const_271;
  wire Const_272;
  wire Const_273;
  wire [2:0] Const_274;
  wire Const_275;
  wire [2:0] Const_276;
  wire Const_277;
  wire [2:0] Const_278;
  wire Const_279;
  wire [2:0] Const_280;
  wire Const_281;
  wire Const_282;
  wire [2:0] Const_283;
  wire Const_284;
  wire Const_285;
  wire Const_286;
  wire Const_287;
  wire Const_288;
  wire Const_289;
  wire Const_290;
  wire Const_291;
  wire Const_292;
  wire Const_293;
  wire Const_294;
  wire Const_295;
  wire Const_296;
  wire Const_297;
  wire Const_298;
  wire Const_299;
  wire Const_300;
  wire Const_301;
  wire Const_302;
  wire Const_303;
  wire Const_304;
  wire Const_305;
  wire Const_306;
  wire Const_307;
  wire Const_308;
  wire Const_309;
  wire Const_310;
  wire Const_311;
  wire Const_312;
  wire Const_313;
  wire Const_314;
  wire Const_315;
  wire Const_316;
  wire Const_317;
  wire Const_318;
  wire Const_319;
  wire Const_320;
  wire Const_321;
  wire Const_322;
  wire Const_323;
  wire Const_324;
  wire Const_325;
  wire Const_326;
  wire Const_327;
  wire Const_328;
  wire [15:0] Const_329;
  wire Const_330;
  wire Const_331;
  wire Const_332;
  wire Const_333;
  wire Const_334;
  wire Const_335;
  wire Const_336;
  wire Const_337;
  wire Const_338;
  wire Const_339;
  wire Const_340;
  wire Const_341;
  wire Const_342;
  wire Const_343;
  wire Const_344;
  wire Const_345;
  wire Const_346;
  wire Const_347;
  wire Const_348;
  wire Const_349;
  wire Const_350;
  wire Const_351;
  wire Const_352;
  wire Const_353;
  wire Const_354;
  wire Const_355;
  wire Const_356;
  wire Const_357;
  wire Const_358;
  wire Const_359;
  wire Const_360;
  wire Const_361;
  wire Const_362;
  wire Const_363;
  wire Const_364;
  wire Const_365;
  wire Const_366;
  wire Const_367;
  wire Const_368;
  wire Const_369;
  wire [3:0] Const_370;
  wire Const_371;
  wire [3:0] Const_372;
  wire Const_373;
  wire [3:0] Const_374;
  wire Const_375;
  wire [3:0] Const_376;
  wire Const_377;
  wire Const_378;
  wire Const_379;
  wire Const_380;
  wire Const_381;
  wire Const_382;
  wire Const_383;
  wire Const_384;
  wire [3:0] Const_385;
  wire Const_386;
  wire [3:0] Const_387;
  wire Const_388;
  wire [3:0] Const_389;
  wire Const_390;
  wire [3:0] Const_391;
  wire Const_392;
  wire Const_393;
  wire [3:0] Const_394;
  wire Const_395;
  wire Const_396;
  wire Const_397;
  wire Const_398;
  wire [3:0] Const_399;
  wire Const_400;
  wire [3:0] Const_401;
  wire Const_402;
  wire [3:0] Const_403;
  wire Const_404;
  wire [3:0] Const_405;
  wire Const_406;
  wire Const_407;
  wire Const_408;
  wire Const_409;
  wire Const_410;
  wire Const_411;
  wire Const_412;
  wire Const_413;
  wire Const_414;
  wire [3:0] Const_415;
  wire Const_416;
  wire [3:0] Const_417;
  wire Const_418;
  wire [3:0] Const_419;
  wire Const_420;
  wire [3:0] Const_421;
  wire Const_422;
  wire [3:0] Const_423;
  wire Const_424;
  wire Const_425;
  wire Const_426;
  wire Const_427;
  wire Const_428;
  wire Const_429;
  wire Const_430;
  wire Const_431;
  wire Const_432;
  wire Const_433;
  wire Const_434;
  wire Const_435;
  wire Const_436;
  wire Const_437;
  wire Const_438;
  wire Const_439;
  wire Const_440;
  wire Const_441;
  wire Const_442;
  wire Const_443;
  wire Const_444;
  wire Const_445;
  wire Const_446;
  wire Const_447;
  wire Const_448;
  wire Const_449;
  wire Const_450;
  wire Const_451;
  wire Const_452;
  wire Const_453;
  wire Const_454;
  wire Const_455;
  wire Const_456;
  wire Const_457;
  wire Const_458;
  wire Const_459;
  wire Const_460;
  wire Const_461;
  wire Const_462;
  wire Const_463;
  wire Const_464;
  wire Const_465;
  wire Const_466;
  wire Const_467;
  wire Const_468;
  wire Const_469;
  wire Const_470;
  wire Const_471;
  wire Const_472;
  wire Const_473;
  wire Const_474;
  wire [63:0] Const_475;
  wire Const_476;
  wire Const_477;
  wire Const_478;
  wire Const_479;
  wire Const_480;
  wire Const_481;
  wire Const_482;
  wire Const_483;
  wire Const_484;
  wire Const_485;
  wire Const_486;
  wire Const_487;
  wire Const_488;
  wire Const_489;
  wire Const_490;
  wire Const_491;
  wire Const_492;
  wire Const_493;
  wire Const_494;
  wire Const_495;
  wire Const_496;
  wire Const_497;
  wire Const_498;
  wire Const_499;
  wire Const_500;
  wire Const_501;
  wire Const_502;
  wire Const_503;
  wire Const_504;
  wire Const_505;
  wire Const_506;
  wire Const_507;
  wire Const_508;
  wire Const_509;
  wire Const_510;
  wire Const_511;
  wire Const_512;
  wire Const_513;
  wire [3:0] Const_514;
  wire Const_515;
  wire [3:0] Const_516;
  wire Const_517;
  wire Const_518;
  wire Const_519;
  wire Const_520;
  wire Const_521;
  wire Const_522;
  wire Const_523;
  wire Const_524;
  wire Const_525;
  wire Const_526;
  wire Const_527;
  wire Const_528;
  wire Const_529;
  wire Const_530;
  wire Const_531;
  wire Const_532;
  wire Const_533;
  wire Const_534;
  wire Const_535;
  wire Const_536;
  wire Const_537;
  wire Const_538;
  wire Const_539;
  wire Const_540;
  wire Const_541;
  wire Const_542;
  wire Const_543;
  wire Const_544;
  wire Const_545;
  wire Const_546;
  wire Const_547;
  wire Const_548;
  wire Const_549;
  wire Const_550;
  wire Const_551;
  wire Const_552;
  wire Const_553;
  wire Const_554;
  wire Const_555;
  wire Const_556;
  wire Const_557;
  wire Const_558;
  wire Const_559;
  wire Const_560;
  wire Const_561;
  wire Const_562;
  wire Const_563;
  wire Const_564;
  wire Const_565;
  wire Const_566;
  wire Const_567;
  wire Const_568;
  wire Const_569;
  wire Const_570;
  wire Const_571;
  wire Const_572;
  wire Const_573;
  wire Const_574;
  wire Const_575;
  wire Const_576;
  wire Const_577;
  wire Const_578;
  wire Const_579;
  wire [7:0] Const_580;
  wire Const_581;
  wire [7:0] Const_582;
  wire Const_583;
  wire [7:0] Const_584;
  wire Const_585;
  wire [7:0] Const_586;
  wire Const_587;
  wire Const_588;
  wire Const_589;
  wire Const_590;
  wire [7:0] Const_591;
  wire Const_592;
  wire Const_593;
  wire Const_594;
  wire Const_595;
  wire Const_596;
  wire Const_597;
  wire Const_598;
  wire Const_599;
  wire Const_600;
  wire Const_601;
  wire Const_602;
  wire Const_603;
  wire [7:0] Const_604;
  wire Const_605;
  wire [7:0] Const_606;
  wire Const_607;
  wire [7:0] Const_608;
  wire Const_609;
  wire Const_610;
  wire Const_611;
  wire Const_612;
  wire Const_613;
  wire Const_614;
  wire Const_615;
  wire Const_616;
  wire Const_617;
  wire Const_618;
  wire Const_619;
  wire Const_620;
  wire Const_621;
  wire Const_622;
  wire Const_623;
  wire Const_624;
  wire Const_625;
  wire Const_626;
  wire Const_627;
  wire Const_628;
  wire Const_629;
  wire Const_630;
  wire Const_631;
  wire Const_632;
  wire Const_633;
  wire Const_634;
  wire Const_635;
  wire Const_636;
  wire Const_637;
  wire Const_638;
  wire Const_639;
  wire Const_640;
  wire Const_641;
  wire Const_642;
  wire Const_643;
  wire Const_644;
  wire Const_645;
  wire Const_646;
  wire Const_647;
  wire Const_648;
  wire Const_649;
  wire Const_650;
  wire Const_651;
  wire Const_652;
  wire Const_653;
  wire Const_654;
  wire Const_655;
  wire Const_656;
  wire Const_657;
  wire Const_658;
  wire Const_659;
  wire Const_660;
  wire Const_661;
  wire Const_662;
  wire Const_663;
  wire Const_664;
  wire Const_665;
  wire Const_666;
  wire Const_667;
  wire Const_668;
  wire Const_669;
  wire Const_670;
  wire Const_671;
  wire Const_672;
  wire Const_673;
  wire Const_674;
  wire Const_675;
  wire Const_676;
  wire Const_677;
  wire Const_678;
  wire Const_679;
  wire Const_680;
  wire Const_681;
  wire Const_682;
  wire Const_683;
  wire Const_684;
  wire Const_685;
  wire Const_686;
  wire Const_687;
  wire Const_688;
  wire Const_689;
  wire Const_690;
  wire Const_691;
  wire Const_692;
  wire Const_693;
  wire Const_694;
  wire Const_695;
  wire [2:0] Const_696;
  wire [2:0] Const_697;
  wire [2:0] Const_698;
  wire [2:0] Const_699;
  wire [2:0] Const_700;
  wire [2:0] Const_701;
  wire [3:0] Const_702;
  wire [3:0] Const_703;
  wire [3:0] Const_704;
  wire [3:0] Const_705;
  wire [3:0] Const_706;
  wire [3:0] Const_707;
  wire [3:0] Const_708;
  wire [63:0] Const_709;
  wire Const_710;
  wire [3:0] Const_711;
  wire [4:0] Const_712;
  wire [4:0] Const_713;
  wire [3:0] Const_714;
  wire [3:0] Const_715;
  wire [3:0] Const_716;
  wire [7:0] Const_717;
  wire [7:0] Const_718;
  wire [7:0] Const_719;
  wire [7:0] Const_720;
  wire [7:0] Const_721;
  wire [7:0] Const_722;
  wire [7:0] Const_723;
  wire [3:0] Const_724;
  wire [7:0] Const_725;
  wire [3:0] Const_726;
  wire [31:0] Const_727;
  wire [3:0] Const_728;
  wire [31:0] Const_729;
  wire [3:0] Const_730;
  wire [7:0] Const_731;
  wire [7:0] Const_732;
  wire [7:0] Const_733;
  wire [7:0] Const_734;
  wire [7:0] Const_735;
  wire [7:0] Const_736;
  wire [7:0] Const_737;
  wire [7:0] Const_738;
  wire [15:0] Const_739;
  wire [15:0] Const_740;
  wire [15:0] Const_741;
  wire [15:0] Const_742;
  wire [15:0] Const_743;
  wire [15:0] Const_744;
  wire [15:0] Const_745;
  wire [15:0] Const_746;
  wire [15:0] Const_747;
  wire [15:0] Const_748;
  wire [2:0] Const_749;
  wire [15:0] Const_750;
  wire Const_751;
  wire Const_752;
  wire [15:0] Const_753;
  wire [15:0] Const_754;
  wire [15:0] Const_755;
  wire [15:0] Const_756;
  wire [3:0] Const_757;
  wire [3:0] Const_758;
  wire [3:0] Const_759;
  wire [63:0] Const_760;
  wire Const_761;
  wire Const_762;
  wire [31:0] Const_763;
  wire Const_764;
  wire Const_765;
  wire [7:0] Const_766;
  wire Const_767;
  wire Const_768;
  wire [23:0] Const_769;
  wire Const_770;
  wire Const_771;
  wire [15:0] Const_772;
  wire Const_773;
  wire Const_774;
  wire [7:0] Const_775;
  wire Const_776;
  wire Const_777;
  wire Const_778;
  wire Const_779;
  wire Const_780;
  wire [23:0] Const_781;
  wire Const_782;
  wire Const_783;
  wire [15:0] Const_784;
  wire Const_785;
  wire Const_786;
  wire [7:0] Const_787;
  wire Const_788;
  wire Const_789;
  wire [15:0] Const_790;
  wire Const_791;
  wire Const_792;
  wire [3:0] Const_793;
  wire Const_794;
  wire Const_795;
  wire Const_796;
  wire Const_797;
  wire [7:0] Const_798;
  wire Const_799;
  wire Const_800;
  wire [63:0] Const_801;
  wire Const_802;
  wire Const_803;
  wire [3:0] Const_804;
  wire Const_805;
  wire Const_806;
  wire [3:0] Const_807;
  wire Const_808;
  wire Const_809;
  wire [3:0] Const_810;
  wire Const_811;
  wire Const_812;
  wire [3:0] Const_813;
  wire Const_814;
  wire Const_815;
  wire Const_816;
  wire Const_817;
  wire Const_818;
  wire Const_819;
  wire [15:0] Const_820;
  wire Const_821;
  wire Const_822;
  wire [31:0] Const_823;
  wire Const_824;
  wire Const_825;
  wire Const_826;
  wire Const_827;
  wire [3:0] Const_828;
  wire Const_829;
  wire Const_830;
  wire [15:0] Const_831;
  wire Const_832;
  wire Const_833;
  wire [15:0] Const_834;
  wire Const_835;
  wire Const_836;
  wire [6:0] Const_837;
  wire Const_838;
  wire Const_839;
  wire [1:0] Const_840;
  wire Const_841;
  wire Const_842;
  wire [6:0] Const_843;
  wire Const_844;
  wire Const_845;
  wire [1:0] Const_846;
  wire Const_847;
  wire Const_848;
  wire [6:0] Const_849;
  wire Const_850;
  wire Const_851;
  wire [2:0] Const_852;
  wire Const_853;
  wire Const_854;
  wire [6:0] Const_855;
  wire Const_856;
  wire Const_857;
  wire [2:0] Const_858;
  wire Const_859;
  wire Const_860;
  wire [6:0] Const_861;
  wire Const_862;
  wire Const_863;
  wire [3:0] Const_864;
  wire Const_865;
  wire Const_866;
  wire [6:0] Const_867;
  wire Const_868;
  wire Const_869;
  wire [3:0] Const_870;
  wire Const_871;
  wire Const_872;
  wire [6:0] Const_873;
  wire Const_874;
  wire Const_875;
  wire [4:0] Const_876;
  wire Const_877;
  wire Const_878;
  wire [6:0] Const_879;
  wire Const_880;
  wire Const_881;
  wire [4:0] Const_882;
  wire Const_883;
  wire Const_884;
  wire [1:0] Const_885;
  wire Const_886;
  wire Const_887;
  wire [1:0] Const_888;
  wire Const_889;
  wire Const_890;
  wire [1:0] Const_891;
  wire Const_892;
  wire Const_893;
  wire [16:0] Const_894;
  wire Const_895;
  wire Const_896;
  wire [16:0] Const_897;
  wire Const_898;
  wire Const_899;
  wire [16:0] Const_900;
  wire Const_901;
  wire Const_902;
  wire [1:0] Const_903;
  wire Const_904;
  wire Const_905;
  wire [16:0] Const_906;
  wire Const_907;
  wire Const_908;
  wire [1:0] Const_909;
  wire Const_910;
  wire Const_911;
  wire [16:0] Const_912;
  wire Const_913;
  wire Const_914;
  wire [1:0] Const_915;
  wire Const_916;
  wire Const_917;
  wire [1:0] Const_918;
  wire Const_919;
  wire Const_920;
  wire [1:0] Const_921;
  wire Const_922;
  wire Const_923;
  wire [16:0] Const_924;
  wire Const_925;
  wire Const_926;
  wire [1:0] Const_927;
  wire Const_928;
  wire Const_929;
  wire [16:0] Const_930;
  wire Const_931;
  wire Const_932;
  wire [15:0] Const_933;
  wire Const_934;
  wire Const_935;
  wire [15:0] Const_936;
  wire Const_937;
  wire Const_938;
  wire [7:0] Const_939;
  wire Const_940;
  wire Const_941;
  wire Const_942;
  wire Const_943;
  wire [15:0] Const_944;
  wire Const_945;
  wire Const_946;
  wire [15:0] Const_947;
  wire Const_948;
  wire Const_949;
  wire [5:0] Const_950;
  wire Const_951;
  wire Const_952;
  wire [15:0] Const_953;
  wire Const_954;
  wire Const_955;
  wire [5:0] Const_956;
  wire Const_957;
  wire Const_958;
  wire [7:0] Const_959;
  wire Const_960;
  wire Const_961;
  wire [7:0] Const_962;
  wire [4:0] Const_963;
  wire [4:0] Const_964;
  wire [7:0] Const_965;
  wire [14:0] Const_966;
  wire [31:0] Const_967;
  wire [14:0] Const_968;
  wire [14:0] Const_969;
  wire [14:0] Const_970;
  wire [31:0] Const_971;
  wire Const_972;
  wire Const_973;
  wire Const_974;
  wire Const_975;
  wire [4:0] Const_976;
  wire [4:0] Const_977;
  wire Const_978;
  wire [23:0] Const_979;
  wire [23:0] Const_980;
  wire Const_981;
  wire [31:0] Const_982;
  wire [31:0] Const_983;
  wire Const_984;
  wire [23:0] Const_985;
  wire [23:0] Const_986;
  wire Const_987;
  wire [15:0] Const_988;
  wire [15:0] Const_989;
  wire Const_990;
  wire [7:0] Const_991;
  wire [7:0] Const_992;
  wire Const_993;
  wire [31:0] Const_994;
  wire [31:0] Const_995;
  wire Const_996;
  wire Const_997;
  wire Const_998;
  wire [4:0] Const_999;
  wire Const_1000;
  wire [63:0] Const_1001;
  wire [63:0] Const_1002;
  wire Const_1003;
  wire Const_1004;
  wire Const_1005;
  wire Const_1006;
  wire [7:0] Const_1007;
  wire [7:0] Const_1008;
  wire Const_1009;
  wire Const_1010;
  wire [7:0] Const_1011;
  wire [7:0] Const_1012;
  wire Const_1013;
  wire Const_1014;
  wire [7:0] Const_1015;
  wire [7:0] Const_1016;
  wire Const_1017;
  wire Const_1018;
  wire [7:0] Const_1019;
  wire [7:0] Const_1020;
  wire Const_1021;
  wire Const_1022;
  wire [7:0] Const_1023;
  wire [7:0] Const_1024;
  wire Const_1025;
  wire Const_1026;
  wire [7:0] Const_1027;
  wire [7:0] Const_1028;
  wire Const_1029;
  wire Const_1030;
  wire [7:0] Const_1031;
  wire [7:0] Const_1032;
  wire Const_1033;
  wire Const_1034;
  wire [7:0] Const_1035;
  wire [7:0] Const_1036;
  wire Const_1037;
  wire [6:0] Const_1038;
  wire Const_1039;
  wire [6:0] Const_1040;
  wire Const_1041;
  wire [6:0] Const_1042;
  wire Const_1043;
  wire [6:0] Const_1044;
  wire Const_1045;
  wire [6:0] Const_1046;
  wire Const_1047;
  wire Const_1048;
  wire [15:0] Const_1049;
  wire [15:0] Const_1050;
  wire Const_1051;
  wire Const_1052;
  wire [15:0] Const_1053;
  wire [15:0] Const_1054;
  wire Const_1055;
  wire Const_1056;
  wire [6:0] Const_1057;
  wire Const_1058;
  wire [6:0] Const_1059;
  wire Const_1060;
  wire [6:0] Const_1061;
  wire Const_1062;
  wire [15:0] Const_1063;
  wire [15:0] Const_1064;
  wire Const_1065;
  wire Const_1066;
  wire [5:0] Const_1067;
  wire [5:0] Const_1068;
  wire Const_1069;
  wire [14:0] Const_1070;
  wire Const_1071;
  wire [15:0] Const_1072;
  wire Const_1073;
  wire [15:0] Const_1074;
  wire [63:0] Const_1075;
  wire [15:0] Const_1076;
  wire Const_1077;
  wire [15:0] Const_1078;
  wire [31:0] Const_1079;
  wire [15:0] Const_1080;
  wire [5:0] Const_1081;
  wire [14:0] Const_1082;
  wire [15:0] Const_1083;
  wire [15:0] Const_1084;
  wire [7:0] Const_1085;
  wire [16:0] Const_1086;
  wire [16:0] Const_1087;
  wire [16:0] Const_1088;
  wire [16:0] Const_1089;
  wire [16:0] Const_1090;
  wire [16:0] Const_1091;
  wire [16:0] Const_1092;
  wire [16:0] Const_1093;
  wire [16:0] Const_1094;
  wire [16:0] Const_1095;
  wire Const_1096;
  wire [15:0] Const_1097;
  wire Const_1098;
  wire [15:0] Const_1099;
  wire [15:0] Const_1100;
  wire [15:0] Const_1101;
  wire Const_1102;
  wire Const_1103;
  wire Const_1104;
  wire Const_1105;
  wire [15:0] Const_1106;
  wire Const_1107;
  wire [15:0] Const_1108;
  wire Const_1109;
  wire [15:0] Const_1110;
  wire Const_1111;
  wire Const_1112;
  wire Const_1113;
  wire Const_1114;
  wire Const_1115;
  wire Const_1116;
  wire Const_1117;
  input [6142:0] locking_key;
  wire [4656:0] working_key;

  initial begin
    #0 ap_CS_fsm = 60'd1;
  end


  Gsm_LPC_Analysis_bkb
  #(
    .DataWidth(4),
    .AddressRange(256),
    .AddressWidth(8)
  )
  bitoff_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(bitoff_address0),
    .ce0(bitoff_ce0),
    .q0(bitoff_q0),
    .address1(bitoff_address1),
    .ce1(bitoff_ce1),
    .q1(bitoff_q1),
    .address2(bitoff_address2),
    .ce2(bitoff_ce2),
    .q2(bitoff_q2),
    .address3(bitoff_address3),
    .ce3(bitoff_ce3),
    .q3(bitoff_q3)
  );


  Gsm_LPC_Analysis_cud
  #(
    .DataWidth(16),
    .AddressRange(9),
    .AddressWidth(4)
  )
  ACF_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(ACF_address0),
    .ce0(ACF_ce0),
    .we0(ACF_we0),
    .d0(ACF_d0),
    .q0(ACF_q0)
  );


  Gsm_LPC_Analysis_cud
  #(
    .DataWidth(16),
    .AddressRange(9),
    .AddressWidth(4)
  )
  P_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(P_address0),
    .ce0(P_ce0),
    .we0(P_we0),
    .d0(P_d0),
    .q0(P_q0)
  );


  Gsm_LPC_Analysis_cud
  #(
    .DataWidth(16),
    .AddressRange(9),
    .AddressWidth(4)
  )
  K_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(K_address0),
    .ce0(K_ce0),
    .we0(K_we0),
    .d0(K_d0),
    .q0(K_q0)
  );


  Gsm_LPC_Analysis_dEe
  #(
    .DataWidth(64),
    .AddressRange(9),
    .AddressWidth(4)
  )
  L_ACF_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(L_ACF_address0),
    .ce0(L_ACF_ce0),
    .we0(L_ACF_we0),
    .d0(L_ACF_d0),
    .q0(L_ACF_q0),
    .address1(L_ACF_address1),
    .ce1(L_ACF_ce1),
    .we1(L_ACF_we1),
    .d1(L_ACF_d1),
    .q1(L_ACF_q1)
  );


  GSM_mac_muladd_15eOg
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(15),
    .din1_WIDTH(16),
    .din2_WIDTH(16),
    .dout_WIDTH(31)
  )
  GSM_mac_muladd_15eOg_U1
  (
    .din0(grp_fu_4288_p0),
    .din1(s_q0),
    .din2(grp_fu_4288_p2),
    .dout(grp_fu_4288_p3)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U2
  (
    .din0(mul_ln93_fu_4296_p0),
    .din1(mul_ln93_fu_4296_p1),
    .dout(mul_ln93_fu_4296_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U3
  (
    .din0(mul_ln94_fu_4302_p0),
    .din1(mul_ln94_fu_4302_p1),
    .dout(mul_ln94_fu_4302_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U4
  (
    .din0(mul_ln98_fu_4308_p0),
    .din1(mul_ln98_fu_4308_p1),
    .dout(mul_ln98_fu_4308_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U5
  (
    .din0(mul_ln100_fu_4314_p0),
    .din1(mul_ln100_fu_4314_p1),
    .dout(mul_ln100_fu_4314_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U6
  (
    .din0(mul_ln103_fu_4320_p0),
    .din1(mul_ln103_fu_4320_p1),
    .dout(mul_ln103_fu_4320_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U7
  (
    .din0(mul_ln107_fu_4326_p0),
    .din1(mul_ln107_fu_4326_p1),
    .dout(mul_ln107_fu_4326_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U8
  (
    .din0(sl_5_reg_4794),
    .din1(mul_ln116_fu_4332_p1),
    .dout(mul_ln116_fu_4332_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U9
  (
    .din0(mul_ln118_fu_4338_p0),
    .din1(mul_ln118_fu_4338_p1),
    .dout(mul_ln118_fu_4338_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U10
  (
    .din0(mul_ln120_fu_4344_p0),
    .din1(mul_ln120_fu_4344_p1),
    .dout(mul_ln120_fu_4344_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U11
  (
    .din0(mul_ln121_fu_4350_p0),
    .din1(mul_ln121_fu_4350_p1),
    .dout(mul_ln121_fu_4350_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U12
  (
    .din0(mul_ln122_fu_4356_p0),
    .din1(mul_ln122_fu_4356_p1),
    .dout(mul_ln122_fu_4356_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U13
  (
    .din0(mul_ln123_fu_4362_p0),
    .din1(mul_ln123_fu_4362_p1),
    .dout(mul_ln123_fu_4362_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U14
  (
    .din0(mul_ln124_fu_4368_p0),
    .din1(mul_ln124_fu_4368_p1),
    .dout(mul_ln124_fu_4368_p2)
  );


  GSM_am_addmul_16sg8j
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(16),
    .dout_WIDTH(33)
  )
  GSM_am_addmul_16sg8j_U15
  (
    .din0(sl_1_reg_4732),
    .din1(sl_3_reg_4760),
    .din2(sl_2_reg_4754),
    .dout(grp_fu_4374_p3)
  );


  GSM_am_addmul_16sg8j
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(16),
    .dout_WIDTH(33)
  )
  GSM_am_addmul_16sg8j_U16
  (
    .din0(sl_5_reg_4794),
    .din1(s_q0),
    .din2(s_q1),
    .dout(grp_fu_4382_p3)
  );


  GSM_mac_muladd_16hbi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(32),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16hbi_U17
  (
    .din0(grp_fu_4390_p0),
    .din1(grp_fu_4390_p1),
    .din2(mul_ln100_reg_4861),
    .dout(grp_fu_4390_p3)
  );


  GSM_mac_muladd_16ibs
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(33),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16ibs_U18
  (
    .din0(grp_fu_4397_p0),
    .din1(grp_fu_4397_p1),
    .din2(grp_fu_4447_p3),
    .dout(grp_fu_4397_p3)
  );


  GSM_mac_muladd_16hbi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(32),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16hbi_U19
  (
    .din0(grp_fu_4403_p0),
    .din1(grp_fu_4403_p1),
    .din2(mul_ln98_reg_4844),
    .dout(grp_fu_4403_p3)
  );


  GSM_mac_muladd_16hbi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(32),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16hbi_U20
  (
    .din0(grp_fu_4410_p0),
    .din1(grp_fu_4410_p1),
    .din2(mul_ln118_reg_4917),
    .dout(grp_fu_4410_p3)
  );


  GSM_mac_muladd_16hbi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(32),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16hbi_U21
  (
    .din0(grp_fu_4416_p0),
    .din1(grp_fu_4416_p1),
    .din2(mul_ln103_reg_4866),
    .dout(grp_fu_4416_p3)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U22
  (
    .din0(mul_ln109_fu_4422_p0),
    .din1(mul_ln109_fu_4422_p1),
    .dout(mul_ln109_fu_4422_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U23
  (
    .din0(mul_ln111_fu_4426_p0),
    .din1(mul_ln111_fu_4426_p1),
    .dout(mul_ln111_fu_4426_p2)
  );


  GSM_mac_muladd_16hbi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(32),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16hbi_U24
  (
    .din0(grp_fu_4430_p0),
    .din1(grp_fu_4430_p1),
    .din2(mul_ln107_reg_4880),
    .dout(grp_fu_4430_p3)
  );


  GSM_mac_muladd_16ibs
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(33),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16ibs_U25
  (
    .din0(grp_fu_4437_p0),
    .din1(grp_fu_4437_p1),
    .din2(grp_fu_4473_p3),
    .dout(grp_fu_4437_p3)
  );


  GSM_mac_muladd_16ibs
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(33),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16ibs_U26
  (
    .din0(grp_fu_4442_p0),
    .din1(grp_fu_4442_p1),
    .din2(grp_fu_4481_p3),
    .dout(grp_fu_4442_p3)
  );


  GSM_mac_muladd_16hbi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(32),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16hbi_U27
  (
    .din0(grp_fu_4447_p0),
    .din1(grp_fu_4447_p1),
    .din2(mul_ln93_reg_4826),
    .dout(grp_fu_4447_p3)
  );


  GSM_ama_addmuladdjbC
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(16),
    .din3_WIDTH(33),
    .dout_WIDTH(34)
  )
  GSM_ama_addmuladdjbC_U28
  (
    .din0(grp_fu_4456_p0),
    .din1(grp_fu_4456_p1),
    .din2(sl_4_reg_4788),
    .din3(mul_ln127_2_reg_4952),
    .dout(grp_fu_4456_p4)
  );


  GSM_mac_muladd_16hbi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(32),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16hbi_U29
  (
    .din0(grp_fu_4465_p0),
    .din1(grp_fu_4465_p1),
    .din2(mul_ln120_reg_4922),
    .dout(grp_fu_4465_p3)
  );


  GSM_mac_muladd_16hbi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(32),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16hbi_U30
  (
    .din0(grp_fu_4473_p0),
    .din1(grp_fu_4473_p1),
    .din2(mul_ln121_reg_4927),
    .dout(grp_fu_4473_p3)
  );


  GSM_mac_muladd_16hbi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(32),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16hbi_U31
  (
    .din0(grp_fu_4481_p0),
    .din1(grp_fu_4481_p1),
    .din2(mul_ln122_reg_4932),
    .dout(grp_fu_4481_p3)
  );


  GSM_mac_muladd_16hbi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(32),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16hbi_U32
  (
    .din0(grp_fu_4489_p0),
    .din1(grp_fu_4489_p1),
    .din2(mul_ln123_reg_4937),
    .dout(grp_fu_4489_p3)
  );


  GSM_mac_muladd_16hbi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(32),
    .dout_WIDTH(33)
  )
  GSM_mac_muladd_16hbi_U33
  (
    .din0(grp_fu_4497_p0),
    .din1(grp_fu_4497_p1),
    .din2(mul_ln124_reg_4942),
    .dout(grp_fu_4497_p3)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U34
  (
    .din0(mul_ln133_fu_4504_p0),
    .din1(mul_ln133_fu_4504_p1),
    .dout(mul_ln133_fu_4504_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U35
  (
    .din0(s_q1),
    .din1(mul_ln141_fu_4509_p1),
    .dout(mul_ln141_fu_4509_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U36
  (
    .din0(s_q0),
    .din1(mul_ln142_fu_4515_p1),
    .dout(mul_ln142_fu_4515_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U37
  (
    .din0(mul_ln140_fu_4521_p0),
    .din1(mul_ln140_fu_4521_p1),
    .dout(mul_ln140_fu_4521_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U38
  (
    .din0(s_q1),
    .din1(mul_ln143_fu_4525_p1),
    .dout(mul_ln143_fu_4525_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U39
  (
    .din0(s_q0),
    .din1(mul_ln144_fu_4530_p1),
    .dout(mul_ln144_fu_4530_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U40
  (
    .din0(s_q1),
    .din1(mul_ln145_fu_4535_p1),
    .dout(mul_ln145_fu_4535_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U41
  (
    .din0(s_q0),
    .din1(mul_ln146_fu_4540_p1),
    .dout(mul_ln146_fu_4540_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U42
  (
    .din0(s_q1),
    .din1(mul_ln147_fu_4545_p1),
    .dout(mul_ln147_fu_4545_p2)
  );


  GSM_mul_mul_16s_1fYi
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mul_mul_16s_1fYi_U43
  (
    .din0(s_q0),
    .din1(mul_ln148_fu_4550_p1),
    .dout(mul_ln148_fu_4550_p2)
  );


  GSM_mac_muladd_16kbM
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mac_muladd_16kbM_U44
  (
    .din0(temp_3_reg_5366),
    .din1(select_ln213_reg_5434),
    .din2(grp_fu_4555_p2),
    .dout(grp_fu_4555_p3)
  );


  GSM_mac_muladd_16kbM
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mac_muladd_16kbM_U45
  (
    .din0(K_q0),
    .din1(grp_fu_4564_p1),
    .din2(grp_fu_4564_p2),
    .dout(grp_fu_4564_p3)
  );


  GSM_mac_muladd_16kbM
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(16),
    .din2_WIDTH(16),
    .dout_WIDTH(32)
  )
  GSM_mac_muladd_16kbM_U46
  (
    .din0(grp_fu_4572_p0),
    .din1(P_q0),
    .din2(grp_fu_4572_p2),
    .dout(grp_fu_4572_p3)
  );


  GSM_mul_mul_16s_1lbW
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(15),
    .dout_WIDTH(31)
  )
  GSM_mul_mul_16s_1lbW_U47
  (
    .din0(LARc_q1),
    .din1(mul_ln50_fu_4580_p1),
    .dout(mul_ln50_fu_4580_p2)
  );


  GSM_mul_mul_16s_1lbW
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(15),
    .dout_WIDTH(31)
  )
  GSM_mul_mul_16s_1lbW_U48
  (
    .din0(LARc_q1),
    .din1(mul_ln50_1_fu_4587_p1),
    .dout(mul_ln50_1_fu_4587_p2)
  );


  GSM_mul_mul_16s_1lbW
  #(
    .ID(1),
    .NUM_STAGE(1),
    .din0_WIDTH(16),
    .din1_WIDTH(15),
    .dout_WIDTH(31)
  )
  GSM_mul_mul_16s_1lbW_U49
  (
    .din0(LARc_q0),
    .din1(mul_ln50_2_fu_4594_p1),
    .dout(mul_ln50_2_fu_4594_p2)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end

  assign Const_16 = (1'd0 ^ working_key[21]);
  assign Const_17 = (1'd1 ^ working_key[22]);
  assign Const_18 = (1'd1 ^ working_key[23]);
  assign Const_19 = (1'd1 ^ working_key[24]);
  assign Const_20 = (1'd0 ^ working_key[25]);
  assign Const_21 = (1'd1 ^ working_key[26]);
  assign Const_22 = (1'd0 ^ working_key[27]);
  assign Const_23 = (1'd0 ^ working_key[28]);

  always @(posedge ap_clk) begin
    if(((icmp_ln147_fu_2573_p2 == Const_16) & (icmp_ln204_fu_2555_p2 == Const_17) & (Const_18 == ap_CS_fsm_state43) ^ working_key[29]) == 1'b0) begin
      L_num_0_i_i_reg_1006 <= sext_ln138_fu_2561_p1;
    end else if((icmp_ln150_fu_2589_p2 == Const_19) & (icmp_ln147_reg_5407 == Const_20) & (icmp_ln204_reg_5387 == Const_21) & (icmp_ln178_reg_5248 == Const_22) & (Const_23 == ap_CS_fsm_state44)) begin
      L_num_0_i_i_reg_1006 <= L_num_3_fu_2611_p3;
    end 
  end

  assign Const_24 = (1'd0 ^ working_key[30]);
  assign Const_25 = (1'd1 ^ working_key[31]);
  assign Const_26 = (1'd1 ^ working_key[32]);
  assign Const_27 = (16'd13641 ^ working_key[48:33]);
  assign Const_28 = (1'd1 ^ working_key[49]);
  assign Const_29 = (1'd0 ^ working_key[50]);
  assign Const_30 = (1'd1 ^ working_key[51]);
  assign Const_31 = (1'd1 ^ working_key[52]);
  assign Const_32 = (1'd0 ^ working_key[53]);

  always @(posedge ap_clk) begin
    if(((icmp_ln147_fu_2573_p2 == Const_24) & (icmp_ln204_fu_2555_p2 == Const_25) & (Const_26 == ap_CS_fsm_state43) ^ working_key[54]) == 1'b1) begin
      div_0_i_i_reg_1015 <= Const_27;
    end else if((icmp_ln150_fu_2589_p2 == Const_28) & (icmp_ln147_reg_5407 == Const_29) & (icmp_ln204_reg_5387 == Const_30) & (icmp_ln178_reg_5248 == Const_31) & (Const_32 == ap_CS_fsm_state44)) begin
      div_0_i_i_reg_1015 <= div_fu_2629_p3;
    end 
  end

  assign Const_33 = (1'd0 ^ working_key[55]);
  assign Const_34 = (1'd1 ^ working_key[56]);

  always @(posedge ap_clk) begin
    if(((Const_33 == ap_CS_fsm_state28) ^ working_key[57]) == 1'b0) begin
      empty_57_reg_884 <= add_ln140_reg_5156;
    end else if(Const_34 == ap_CS_fsm_state19) begin
      empty_57_reg_884 <= add_ln126_reg_5029;
    end 
  end

  assign Const_35 = (1'd1 ^ working_key[58]);
  assign Const_36 = (1'd0 ^ working_key[59]);
  assign Const_37 = (4'd6 ^ working_key[63:60]);

  always @(posedge ap_clk) begin
    if(((Const_35 == ap_CS_fsm_state36) ^ working_key[64]) == 1'b0) begin
      i_1_i_reg_928 <= i_reg_5300;
    end else if(Const_36 == ap_CS_fsm_state34) begin
      i_1_i_reg_928 <= Const_37;
    end 
  end

  assign Const_38 = (1'd1 ^ working_key[65]);
  assign Const_39 = (1'd0 ^ working_key[66]);
  assign Const_40 = (4'd5 ^ working_key[70:67]);
  assign Const_41 = (1'd1 ^ working_key[71]);

  always @(posedge ap_clk) begin
    if(((icmp_ln186_fu_2443_p2 == Const_38) & (Const_39 == ap_CS_fsm_state35) ^ working_key[72]) == 1'b0) begin
      i_2_i_reg_939 <= Const_40;
    end else if(Const_41 == ap_CS_fsm_state38) begin
      i_2_i_reg_939 <= i_1_reg_5328;
    end 
  end

  assign Const_42 = (1'd1 ^ working_key[73]);
  assign Const_43 = (1'd0 ^ working_key[74]);
  assign Const_44 = (4'd10 ^ working_key[78:75]);
  assign Const_45 = (1'd0 ^ working_key[79]);

  always @(posedge ap_clk) begin
    if(((icmp_ln192_fu_2480_p2 == Const_42) & (Const_43 == ap_CS_fsm_state37) ^ working_key[80]) == 1'b1) begin
      i_3_i_reg_950 <= Const_44;
    end else if(Const_45 == ap_CS_fsm_state40) begin
      i_3_i_reg_950 <= i_2_reg_5336;
    end 
  end

  assign Const_46 = (1'd1 ^ working_key[81]);
  assign Const_47 = (1'd0 ^ working_key[82]);
  assign Const_48 = (32'd1431644927 ^ working_key[114:83]);
  assign Const_49 = (1'd0 ^ working_key[115]);
  assign Const_50 = (1'd1 ^ working_key[116]);

  always @(posedge ap_clk) begin
    if(((icmp_ln194_fu_2497_p2 == Const_46) & (Const_47 == ap_CS_fsm_state39) ^ working_key[117]) == 1'b0) begin
      i_3_reg_973 <= Const_48;
    end else if((icmp_ln223_fu_2788_p2 == Const_49) & (Const_50 == ap_CS_fsm_state47)) begin
      i_3_reg_973 <= n_1_fu_2809_p2;
    end 
  end

  assign Const_51 = (1'd1 ^ working_key[118]);
  assign Const_52 = (1'd1 ^ working_key[119]);
  assign Const_53 = (32'd1286253216 ^ working_key[151:120]);
  assign Const_54 = (1'd0 ^ working_key[152]);
  assign Const_55 = (1'd1 ^ working_key[153]);

  always @(posedge ap_clk) begin
    if(((icmp_ln194_fu_2497_p2 == Const_51) & (Const_52 == ap_CS_fsm_state39) ^ working_key[154]) == 1'b0) begin
      indvars_iv142_reg_961 <= Const_53;
    end else if((icmp_ln223_fu_2788_p2 == Const_54) & (Const_55 == ap_CS_fsm_state47)) begin
      indvars_iv142_reg_961 <= add_ln199_2_fu_2815_p2;
    end 
  end

  assign Const_56 = (1'd0 ^ working_key[155]);
  assign Const_57 = (1'd1 ^ working_key[156]);
  assign Const_58 = (1'd0 ^ working_key[157]);
  assign Const_59 = (4'd5 ^ working_key[161:158]);
  assign Const_60 = (1'd0 ^ working_key[162]);
  assign Const_61 = (1'd0 ^ working_key[163]);
  assign Const_62 = (1'd1 ^ working_key[164]);
  assign Const_63 = (1'd0 ^ working_key[165]);
  assign Const_64 = (1'd1 ^ working_key[166]);

  always @(posedge ap_clk) begin
    if(((icmp_ln147_fu_2573_p2 == Const_56) & (icmp_ln204_fu_2555_p2 == Const_57) & (Const_58 == ap_CS_fsm_state43) ^ working_key[167]) == 1'b0) begin
      k_0_i_i_reg_1026 <= Const_59;
    end else if((icmp_ln150_fu_2589_p2 == Const_60) & (icmp_ln147_reg_5407 == Const_61) & (icmp_ln204_reg_5387 == Const_62) & (icmp_ln178_reg_5248 == Const_63) & (Const_64 == ap_CS_fsm_state44)) begin
      k_0_i_i_reg_1026 <= add_ln150_fu_2583_p2;
    end 
  end

  assign Const_65 = (1'd1 ^ working_key[168]);
  assign Const_66 = (1'd0 ^ working_key[169]);
  assign Const_67 = (1'd1 ^ working_key[170]);
  assign Const_68 = (8'd77 ^ working_key[178:171]);

  always @(posedge ap_clk) begin
    if(((Const_65 == ap_CS_fsm_state3) ^ working_key[179]) == 1'b0) begin
      k_0_i_reg_851 <= k_reg_4621;
    end else if((ap_start == Const_66) & (Const_67 == ap_CS_fsm_state1)) begin
      k_0_i_reg_851 <= Const_68;
    end 
  end

  assign Const_69 = (1'd0 ^ working_key[180]);
  assign Const_70 = (8'd85 ^ working_key[188:181]);
  assign Const_71 = (1'd0 ^ working_key[189]);

  always @(posedge ap_clk) begin
    if(((Const_69 == ap_CS_fsm_state5) ^ working_key[190]) == 1'b0) begin
      k_1_i_reg_862 <= Const_70;
    end else if(Const_71 == ap_CS_fsm_state8) begin
      k_1_i_reg_862 <= k_1_reg_4704;
    end 
  end

  assign Const_72 = (1'd0 ^ working_key[191]);
  assign Const_73 = (1'd0 ^ working_key[192]);
  assign Const_74 = (1'd1 ^ working_key[193]);
  assign Const_75 = (5'd1 ^ working_key[198:194]);

  always @(posedge ap_clk) begin
    if(((tmp_14_fu_1558_p3 == Const_72) & (Const_73 == ap_CS_fsm_state10) ^ working_key[199]) == 1'b1) begin
      k_2_i_reg_873 <= k_2_fu_1571_p2;
    end else if(Const_74 == ap_CS_fsm_state9) begin
      k_2_i_reg_873 <= Const_75;
    end 
  end

  assign Const_76 = (1'd0 ^ working_key[200]);
  assign Const_77 = (1'd1 ^ working_key[201]);
  assign Const_78 = (5'd29 ^ working_key[206:202]);
  assign Const_79 = (1'd0 ^ working_key[207]);

  always @(posedge ap_clk) begin
    if(((icmp_ln135_fu_1848_p2 == Const_76) & (Const_77 == ap_CS_fsm_state20) ^ working_key[208]) == 1'b1) begin
      k_3_i_reg_906 <= Const_78;
    end else if(Const_79 == ap_CS_fsm_state30) begin
      k_3_i_reg_906 <= k_3_reg_5230;
    end 
  end

  assign Const_80 = (1'd1 ^ working_key[209]);
  assign Const_81 = (1'd0 ^ working_key[210]);
  assign Const_82 = (32'd1431644927 ^ working_key[242:211]);

  always @(posedge ap_clk) begin
    if(((Const_80 == ap_CS_fsm_state49) ^ working_key[243]) == 1'b0) begin
      m_0_i_reg_1060 <= m_reg_5486;
    end else if(Const_81 == ap_CS_fsm_state46) begin
      m_0_i_reg_1060 <= Const_82;
    end 
  end

  assign Const_83 = (1'd1 ^ working_key[244]);
  assign Const_84 = (1'd1 ^ working_key[245]);
  assign Const_85 = (1'd0 ^ working_key[246]);
  assign Const_86 = (1'd0 ^ working_key[247]);
  assign Const_87 = (1'd1 ^ working_key[248]);
  assign Const_88 = (1'd1 ^ working_key[249]);
  assign Const_89 = (1'd0 ^ working_key[250]);
  assign Const_90 = (1'd0 ^ working_key[251]);
  assign Const_91 = (16'd43690 ^ working_key[267:252]);

  always @(posedge ap_clk) begin
    if(((icmp_ln150_fu_2589_p2 == Const_83) & (icmp_ln147_reg_5407 == Const_84) & (icmp_ln204_reg_5387 == Const_85) & (icmp_ln178_reg_5248 == Const_86) & (Const_87 == ap_CS_fsm_state44) ^ working_key[268]) == 1'b1) begin
      p_0_i52_i_reg_1037 <= div_0_i_i_reg_1015;
    end else if((icmp_ln147_fu_2573_p2 == Const_88) & (icmp_ln204_fu_2555_p2 == Const_89) & (Const_90 == ap_CS_fsm_state43)) begin
      p_0_i52_i_reg_1037 <= Const_91;
    end 
  end

  assign Const_92 = (1'd0 ^ working_key[269]);
  assign Const_93 = (1'd1 ^ working_key[270]);
  assign Const_94 = (1'd0 ^ working_key[271]);
  assign Const_95 = (1'd1 ^ working_key[272]);
  assign Const_96 = (1'd1 ^ working_key[273]);
  assign Const_97 = (1'd0 ^ working_key[274]);
  assign Const_98 = (1'd0 ^ working_key[275]);
  assign Const_99 = (1'd0 ^ working_key[276]);
  assign Const_100 = (1'd0 ^ working_key[277]);
  assign Const_101 = (1'd0 ^ working_key[278]);
  assign Const_102 = (1'd1 ^ working_key[279]);
  assign Const_103 = (4'd5 ^ working_key[283:280]);

  always @(posedge ap_clk) begin
    if(((Const_92 == ap_CS_fsm_state53) ^ working_key[284]) == 1'b0) begin
      p_0_rec_i16_reg_1082 <= add_ln253_reg_5541;
    end else if((Const_93 == ap_CS_fsm_state44) & ((icmp_ln178_reg_5248 == Const_94) | ((icmp_ln206_fu_2677_p2 == Const_95) & (icmp_ln204_reg_5387 == Const_96) | (icmp_ln215_fu_2657_p2 == Const_97) & (icmp_ln150_fu_2589_p2 == Const_98) & (icmp_ln204_reg_5387 == Const_99) | (icmp_ln215_fu_2657_p2 == Const_100) & (icmp_ln147_reg_5407 == Const_101) & (icmp_ln204_reg_5387 == Const_102)))) begin
      p_0_rec_i16_reg_1082 <= Const_103;
    end 
  end

  assign Const_104 = (1'd0 ^ working_key[285]);
  assign Const_105 = (1'd1 ^ working_key[286]);
  assign Const_106 = (4'd5 ^ working_key[290:287]);
  assign Const_107 = (1'd0 ^ working_key[291]);
  assign Const_108 = (1'd0 ^ working_key[292]);

  always @(posedge ap_clk) begin
    if(((icmp_ln178_fu_2101_p2 == Const_104) & (Const_105 == ap_CS_fsm_state33) ^ working_key[293]) == 1'b1) begin
      p_0_rec_i1_reg_1071 <= Const_106;
    end else if((icmp_ln180_fu_3008_p2 == Const_107) & (Const_108 == ap_CS_fsm_state50)) begin
      p_0_rec_i1_reg_1071 <= add_ln181_fu_3014_p2;
    end 
  end

  assign Const_109 = (1'd1 ^ working_key[294]);
  assign Const_110 = (1'd0 ^ working_key[295]);
  assign Const_111 = (1'd1 ^ working_key[296]);
  assign Const_112 = (8'd53 ^ working_key[304:297]);
  assign Const_113 = (1'd0 ^ working_key[305]);

  always @(posedge ap_clk) begin
    if(((tmp_15_fu_2052_p3 == Const_109) & (icmp_ln72_reg_4683 == Const_110) & (Const_111 == ap_CS_fsm_state29) ^ working_key[306]) == 1'b1) begin
      p_0_rec_i_reg_917 <= Const_112;
    end else if(Const_113 == ap_CS_fsm_state32) begin
      p_0_rec_i_reg_917 <= add_ln159_reg_5243;
    end 
  end

  assign Const_114 = (1'd0 ^ working_key[307]);
  assign Const_115 = (1'd0 ^ working_key[308]);
  assign Const_116 = (4'd5 ^ working_key[312:309]);
  assign Const_117 = (1'd0 ^ working_key[313]);
  assign Const_118 = (1'd1 ^ working_key[314]);

  always @(posedge ap_clk) begin
    if(((icmp_ln194_fu_2497_p2 == Const_114) & (Const_115 == ap_CS_fsm_state39) ^ working_key[315]) == 1'b0) begin
      p_1_rec_i_reg_985 <= Const_116;
    end else if((icmp_ln223_fu_2788_p2 == Const_117) & (Const_118 == ap_CS_fsm_state47)) begin
      p_1_rec_i_reg_985 <= add_ln199_reg_5377;
    end 
  end

  assign Const_119 = (1'd1 ^ working_key[316]);
  assign Const_120 = (1'd0 ^ working_key[317]);
  assign Const_121 = (32'd1607685269 ^ working_key[349:318]);
  assign Const_122 = (1'd0 ^ working_key[350]);
  assign Const_123 = (1'd0 ^ working_key[351]);
  assign Const_124 = (1'd1 ^ working_key[352]);
  assign Const_125 = (1'd1 ^ working_key[353]);

  always @(posedge ap_clk) begin
    if(((icmp_ln204_fu_2555_p2 == Const_119) & (Const_120 == ap_CS_fsm_state43) ^ working_key[354]) == 1'b1) begin
      p_2_rec_i_reg_1049 <= Const_121;
    end else if((icmp_ln204_reg_5387 == Const_122) & (icmp_ln206_fu_2677_p2 == Const_123) & (icmp_ln178_reg_5248 == Const_124) & (Const_125 == ap_CS_fsm_state44)) begin
      p_2_rec_i_reg_1049 <= add_ln207_fu_2683_p2;
    end 
  end

  assign Const_126 = (1'd0 ^ working_key[355]);
  assign Const_127 = (1'd1 ^ working_key[356]);
  assign Const_128 = (1'd0 ^ working_key[357]);

  always @(posedge ap_clk) begin
    if(((Const_126 == ap_CS_fsm_state21) ^ working_key[358]) == 1'b1) begin
      reg_1099 <= s_q1;
    end else if((Const_127 == ap_CS_fsm_state14) | (Const_128 == ap_CS_fsm_state9)) begin
      reg_1099 <= s_q0;
    end 
  end

  assign Const_129 = (1'd0 ^ working_key[359]);
  assign Const_130 = (1'd1 ^ working_key[360]);
  assign Const_131 = (1'd0 ^ working_key[361]);

  always @(posedge ap_clk) begin
    if((((Const_129 == ap_CS_fsm_state23) | (Const_130 == ap_CS_fsm_state21)) ^ working_key[362]) == 1'b1) begin
      reg_1104 <= L_ACF_q1;
    end else if(Const_131 == ap_CS_fsm_state13) begin
      reg_1104 <= L_ACF_q0;
    end 
  end

  assign Const_132 = (1'd0 ^ working_key[363]);
  assign Const_133 = (1'd1 ^ working_key[364]);
  assign Const_134 = (1'd0 ^ working_key[365]);
  assign Const_135 = (1'd1 ^ working_key[366]);

  always @(posedge ap_clk) begin
    if((((Const_132 == ap_CS_fsm_state23) | (Const_133 == ap_CS_fsm_state21)) ^ working_key[367]) == 1'b0) begin
      reg_1109 <= L_ACF_q0;
    end else if((Const_134 == ap_CS_fsm_state15) | (Const_135 == ap_CS_fsm_state13)) begin
      reg_1109 <= L_ACF_q1;
    end 
  end

  assign Const_136 = (1'd1 ^ working_key[368]);
  assign Const_137 = (1'd0 ^ working_key[369]);
  assign Const_138 = (1'd1 ^ working_key[370]);
  assign Const_139 = (16'd21765 ^ working_key[386:371]);

  always @(posedge ap_clk) begin
    if(((Const_136 == ap_CS_fsm_state3) ^ working_key[387]) == 1'b0) begin
      smax_0_i_reg_839 <= select_ln61_fu_1334_p3;
    end else if((ap_start == Const_137) & (Const_138 == ap_CS_fsm_state1)) begin
      smax_0_i_reg_839 <= Const_139;
    end 
  end

  assign Const_140 = (1'd1 ^ working_key[388]);
  assign Const_141 = (1'd0 ^ working_key[389]);
  assign Const_142 = (8'd170 ^ working_key[397:390]);

  always @(posedge ap_clk) begin
    if(((Const_140 == ap_CS_fsm_state28) ^ working_key[398]) == 1'b1) begin
      sp_0_rec_i_reg_894 <= add_ln138_reg_5073;
    end else if(Const_141 == ap_CS_fsm_state19) begin
      sp_0_rec_i_reg_894 <= Const_142;
    end 
  end

  assign Const_143 = (1'd0 ^ working_key[399]);
  assign Const_144 = (1'd0 ^ working_key[400]);
  assign Const_145 = (1'd1 ^ working_key[401]);

  always @(posedge ap_clk) begin
    if(Const_143 == ap_CS_fsm_state42) begin
      if(((tmp_21_fu_2519_p3 == Const_144) ^ working_key[402]) == 1'b0) begin
        temp_24_reg_997 <= P_q0;
      end else if(tmp_21_fu_2519_p3 == Const_145) begin
        temp_24_reg_997 <= zext_ln72_fu_2551_p1;
      end 
    end 
  end

  assign Const_146 = (1'd1 ^ working_key[403]);
  assign Const_147 = (1'd1 ^ working_key[404]);

  always @(posedge ap_clk) begin
    if((icmp_ln223_fu_2788_p2 == Const_146) & (Const_147 == ap_CS_fsm_state47)) begin
      K_addr_1_reg_5481 <= zext_ln225_fu_2793_p1;
      m_reg_5486 <= m_fu_2798_p2;
      zext_ln225_reg_5476[31:0] <= zext_ln225_fu_2793_p1[31:0];
    end 
  end

  assign Const_148 = (1'd1 ^ working_key[405]);

  always @(posedge ap_clk) begin
    if(Const_148 == ap_CS_fsm_state48) begin
      K_load_reg_5506 <= K_q0;
      temp_6_reg_5512 <= temp_6_fu_2845_p3;
      temp_7_reg_5518 <= temp_7_fu_2871_p3;
    end 
  end

  assign Const_149 = (1'd0 ^ working_key[406]);

  always @(posedge ap_clk) begin
    if(Const_149 == ap_CS_fsm_state42) begin
      LARc_addr_2_reg_5361 <= zext_ln206_fu_2514_p1;
      add_ln199_reg_5377 <= add_ln199_fu_2527_p2;
      temp_3_reg_5366 <= P_q0;
    end 
  end

  assign Const_150 = (1'd1 ^ working_key[407]);

  always @(posedge ap_clk) begin
    if(Const_150 == ap_CS_fsm_state51) begin
      LARc_addr_4_reg_5532 <= p_0_rec_i16_cast_fu_3020_p1;
      add_ln253_reg_5541 <= add_ln253_fu_3031_p2;
    end 
  end

  assign Const_151 = (1'd1 ^ working_key[408]);
  assign Const_152 = (1'd1 ^ working_key[409]);

  always @(posedge ap_clk) begin
    if((tmp_15_fu_2052_p3 == Const_151) & (Const_152 == ap_CS_fsm_state29)) begin
      L_ACF_addr_9_reg_5224 <= zext_ln152_fu_2060_p1;
      k_3_reg_5230 <= k_3_fu_2065_p2;
    end 
  end

  assign Const_153 = (1'd0 ^ working_key[410]);

  always @(posedge ap_clk) begin
    if(Const_153 == ap_CS_fsm_state15) begin
      add_ln126_2_reg_4973 <= grp_fu_4410_p3;
      add_ln126_7_reg_4978 <= add_ln126_7_fu_1672_p2;
      add_ln127_reg_4983 <= add_ln127_fu_1699_p2;
      add_ln128_reg_4988 <= add_ln128_fu_1730_p2;
      add_ln129_1_reg_4993 <= grp_fu_4416_p3;
      add_ln129_4_reg_4998 <= grp_fu_4437_p3;
      add_ln130_3_reg_5003 <= grp_fu_4442_p3;
      add_ln131_reg_5008 <= add_ln131_fu_1745_p2;
      add_ln132_1_reg_5013 <= grp_fu_4497_p3;
      mul_ln109_reg_4957 <= mul_ln109_fu_4422_p2;
      mul_ln111_reg_4962 <= mul_ln111_fu_4426_p2;
      mul_ln133_reg_5018 <= mul_ln133_fu_4504_p2;
    end 
  end

  assign Const_154 = (1'd1 ^ working_key[411]);

  always @(posedge ap_clk) begin
    if(Const_154 == ap_CS_fsm_state16) begin
      add_ln126_reg_5029 <= add_ln126_fu_1775_p2;
      add_ln129_reg_5034 <= add_ln129_fu_1794_p2;
      add_ln130_reg_5039 <= add_ln130_fu_1809_p2;
      add_ln132_reg_5044 <= add_ln132_fu_1818_p2;
      add_ln133_reg_5049 <= add_ln133_fu_1827_p2;
    end 
  end

  assign Const_155 = (1'd0 ^ working_key[412]);

  always @(posedge ap_clk) begin
    if(Const_155 == ap_CS_fsm_state20) begin
      add_ln138_reg_5073 <= add_ln138_fu_1854_p2;
      s_addr_10_reg_5065 <= sum17_cast_fu_1843_p1;
      sp_0_rec_i_cast_reg_5060[7:0] <= sp_0_rec_i_cast_fu_1833_p1[7:0];
    end 
  end

  assign Const_156 = (1'd0 ^ working_key[413]);

  always @(posedge ap_clk) begin
    if(Const_156 == ap_CS_fsm_state24) begin
      add_ln140_reg_5156 <= add_ln140_fu_1971_p2;
      add_ln143_1_reg_5161 <= add_ln143_1_fu_1981_p2;
      add_ln144_1_reg_5166 <= add_ln144_1_fu_1990_p2;
      mul_ln145_reg_5171 <= mul_ln145_fu_4535_p2;
      mul_ln146_reg_5176 <= mul_ln146_fu_4540_p2;
    end 
  end

  assign Const_157 = (1'd1 ^ working_key[414]);

  always @(posedge ap_clk) begin
    if(Const_157 == ap_CS_fsm_state23) begin
      add_ln141_reg_5126 <= add_ln141_fu_1919_p2;
      add_ln142_1_reg_5131 <= add_ln142_1_fu_1928_p2;
      mul_ln140_reg_5121 <= mul_ln140_fu_4521_p2;
      mul_ln143_reg_5136 <= mul_ln143_fu_4525_p2;
      mul_ln144_reg_5141 <= mul_ln144_fu_4530_p2;
    end 
  end

  assign Const_158 = (1'd0 ^ working_key[415]);

  always @(posedge ap_clk) begin
    if(Const_158 == ap_CS_fsm_state25) begin
      add_ln145_1_reg_5191 <= add_ln145_1_fu_2007_p2;
      add_ln146_1_reg_5196 <= add_ln146_1_fu_2016_p2;
      mul_ln147_reg_5201 <= mul_ln147_fu_4545_p2;
      mul_ln148_reg_5206 <= mul_ln148_fu_4550_p2;
    end 
  end

  assign Const_159 = (1'd1 ^ working_key[416]);

  always @(posedge ap_clk) begin
    if(Const_159 == ap_CS_fsm_state26) begin
      add_ln147_reg_5211 <= add_ln147_fu_2033_p2;
      add_ln148_reg_5216 <= add_ln148_fu_2042_p2;
    end 
  end

  assign Const_160 = (1'd0 ^ working_key[417]);
  assign Const_161 = (1'd1 ^ working_key[418]);

  always @(posedge ap_clk) begin
    if((icmp_ln72_reg_4683 == Const_160) & (Const_161 == ap_CS_fsm_state31)) begin
      add_ln159_reg_5243 <= add_ln159_fu_2089_p2;
      s_addr_19_reg_5235 <= p_0_rec_i_cast_fu_2078_p1;
    end 
  end

  assign Const_162 = (1'd1 ^ working_key[419]);

  always @(posedge ap_clk) begin
    if(Const_162 == ap_CS_fsm_state4) begin
      and_ln72_reg_4687 <= and_ln72_fu_1495_p2;
      icmp_ln72_reg_4683 <= icmp_ln72_fu_1483_p2;
      sext_ln67_reg_4678 <= sext_ln67_fu_1479_p1;
    end 
  end

  assign Const_163 = (1'd1 ^ working_key[420]);
  assign Const_164 = (1'd1 ^ working_key[421]);

  always @(posedge ap_clk) begin
    if((icmp_ln192_fu_2480_p2 == Const_163) & (Const_164 == ap_CS_fsm_state37)) begin
      i_1_reg_5328 <= i_1_fu_2491_p2;
      zext_ln193_reg_5318[3:0] <= zext_ln193_fu_2486_p1[3:0];
    end 
  end

  assign Const_165 = (1'd1 ^ working_key[422]);

  always @(posedge ap_clk) begin
    if(Const_165 == ap_CS_fsm_state39) begin
      i_2_reg_5336 <= i_2_fu_2503_p2;
    end 
  end

  assign Const_166 = (1'd0 ^ working_key[423]);

  always @(posedge ap_clk) begin
    if(Const_166 == ap_CS_fsm_state35) begin
      i_reg_5300 <= i_fu_2449_p2;
    end 
  end

  assign Const_167 = (1'd0 ^ working_key[424]);
  assign Const_168 = (1'd0 ^ working_key[425]);

  always @(posedge ap_clk) begin
    if((icmp_ln178_fu_2101_p2 == Const_167) & (Const_168 == ap_CS_fsm_state33)) begin
      icmp_ln118_1_reg_5252 <= icmp_ln118_1_fu_2107_p2;
      or_ln118_2_reg_5287 <= or_ln118_2_fu_2361_p2;
      or_ln118_reg_5282 <= or_ln118_fu_2349_p2;
      sel_tmp57_reg_5277 <= sel_tmp57_fu_2321_p2;
    end 
  end

  assign Const_169 = (1'd1 ^ working_key[426]);
  assign Const_170 = (1'd0 ^ working_key[427]);

  always @(posedge ap_clk) begin
    if((icmp_ln58_fu_1126_p2 == Const_169) & (Const_170 == ap_CS_fsm_state2)) begin
      icmp_ln118_reg_4631 <= icmp_ln118_fu_1151_p2;
      icmp_ln123_1_reg_4648 <= icmp_ln123_1_fu_1231_p2;
      icmp_ln123_2_reg_4668 <= icmp_ln123_2_fu_1286_p2;
      icmp_ln123_reg_4642 <= icmp_ln123_fu_1215_p2;
      tmp_1_reg_4637 <= smax_0_i_reg_839[32'd15];
    end 
  end

  assign Const_171 = (1'd0 ^ working_key[428]);
  assign Const_172 = (1'd0 ^ working_key[429]);

  always @(posedge ap_clk) begin
    if((icmp_ln204_fu_2555_p2 == Const_171) & (Const_172 == ap_CS_fsm_state43)) begin
      icmp_ln147_reg_5407 <= icmp_ln147_fu_2573_p2;
      sext_ln139_1_reg_5402 <= sext_ln139_1_fu_2569_p1;
      sext_ln139_reg_5396 <= sext_ln139_fu_2565_p1;
    end 
  end

  assign Const_173 = (1'd0 ^ working_key[430]);

  always @(posedge ap_clk) begin
    if(Const_173 == ap_CS_fsm_state33) begin
      icmp_ln178_reg_5248 <= icmp_ln178_fu_2101_p2;
    end 
  end

  assign Const_174 = (1'd1 ^ working_key[431]);

  always @(posedge ap_clk) begin
    if(Const_174 == ap_CS_fsm_state43) begin
      icmp_ln204_reg_5387 <= icmp_ln204_fu_2555_p2;
    end 
  end

  assign Const_175 = (1'd1 ^ working_key[432]);

  always @(posedge ap_clk) begin
    if(Const_175 == ap_CS_fsm_state55) begin
      icmp_ln40_10_reg_5587 <= icmp_ln40_10_fu_3423_p2;
      icmp_ln40_8_reg_5597 <= icmp_ln40_8_fu_3495_p2;
      tmp_7_reg_5592 <= { { add_ln40_4_fu_3429_p2[15:9] } };
      tmp_8_reg_5602 <= { { add_ln40_5_fu_3501_p2[15:9] } };
    end 
  end

  assign Const_176 = (1'd0 ^ working_key[433]);

  always @(posedge ap_clk) begin
    if(Const_176 == ap_CS_fsm_state57) begin
      icmp_ln40_12_reg_5643 <= icmp_ln40_12_fu_3790_p2;
      temp_16_reg_5653 <= { { mul_ln50_1_fu_4587_p2[30:15] } };
      temp_17_reg_5659 <= { { mul_ln50_2_fu_4594_p2[30:15] } };
      tmp_9_reg_5648 <= { { add_ln40_8_fu_3796_p2[15:9] } };
    end 
  end

  assign Const_177 = (1'd1 ^ working_key[434]);

  always @(posedge ap_clk) begin
    if(Const_177 == ap_CS_fsm_state56) begin
      icmp_ln40_13_reg_5623 <= icmp_ln40_13_fu_3580_p2;
      temp_13_reg_5617 <= { { mul_ln50_fu_4580_p2[30:15] } };
      tmp_s_reg_5628 <= { { add_ln40_9_fu_3586_p2[15:9] } };
    end 
  end

  assign Const_178 = (1'd0 ^ working_key[435]);

  always @(posedge ap_clk) begin
    if(Const_178 == ap_CS_fsm_state58) begin
      icmp_ln40_14_reg_5665 <= icmp_ln40_14_fu_3977_p2;
      icmp_ln40_15_reg_5675 <= icmp_ln40_15_fu_4007_p2;
      tmp_10_reg_5670 <= { { add_ln40_11_fu_3983_p2[15:9] } };
      tmp_11_reg_5680 <= { { add_ln40_12_fu_4013_p2[15:9] } };
    end 
  end

  assign Const_179 = (1'd0 ^ working_key[436]);

  always @(posedge ap_clk) begin
    if(Const_179 == ap_CS_fsm_state54) begin
      icmp_ln40_6_reg_5557 <= icmp_ln40_6_fu_3219_p2;
      icmp_ln40_7_reg_5567 <= icmp_ln40_7_fu_3301_p2;
      tmp_5_reg_5562 <= { { add_ln40_fu_3225_p2[15:9] } };
      tmp_6_reg_5572 <= { { add_ln40_2_fu_3307_p2[15:9] } };
    end 
  end

  assign Const_180 = (1'd0 ^ working_key[437]);

  always @(posedge ap_clk) begin
    if(Const_180 == ap_CS_fsm_state45) begin
      icmp_ln58_1_reg_5451 <= icmp_ln58_1_fu_2689_p2;
      select_ln40_1_reg_5463 <= select_ln40_1_fu_2774_p3;
      sext_ln62_2_reg_5457 <= sext_ln62_2_fu_2703_p1;
    end 
  end

  assign Const_181 = (1'd1 ^ working_key[438]);
  assign Const_182 = (1'd0 ^ working_key[439]);

  always @(posedge ap_clk) begin
    if((Const_181 == and_ln72_reg_4687) & (Const_182 == ap_CS_fsm_state6)) begin
      k_1_reg_4704 <= k_1_fu_1530_p2;
    end 
  end

  assign Const_183 = (1'd1 ^ working_key[440]);

  always @(posedge ap_clk) begin
    if(Const_183 == ap_CS_fsm_state2) begin
      k_reg_4621 <= k_fu_1132_p2;
    end 
  end

  assign Const_184 = (1'd0 ^ working_key[441]);

  always @(posedge ap_clk) begin
    if(Const_184 == ap_CS_fsm_state14) begin
      mul_ln100_reg_4861 <= mul_ln100_fu_4314_p2;
      mul_ln103_reg_4866 <= mul_ln103_fu_4320_p2;
      mul_ln107_reg_4880 <= mul_ln107_fu_4326_p2;
      mul_ln116_reg_4906 <= mul_ln116_fu_4332_p2;
      mul_ln118_reg_4917 <= mul_ln118_fu_4338_p2;
      mul_ln120_reg_4922 <= mul_ln120_fu_4344_p2;
      mul_ln121_reg_4927 <= mul_ln121_fu_4350_p2;
      mul_ln122_reg_4932 <= mul_ln122_fu_4356_p2;
      mul_ln123_reg_4937 <= mul_ln123_fu_4362_p2;
      mul_ln124_reg_4942 <= mul_ln124_fu_4368_p2;
      mul_ln127_2_reg_4952 <= grp_fu_4382_p3;
      mul_ln127_reg_4947 <= grp_fu_4374_p3;
      mul_ln93_reg_4826 <= mul_ln93_fu_4296_p2;
      mul_ln94_reg_4831 <= mul_ln94_fu_4302_p2;
      mul_ln98_reg_4844 <= mul_ln98_fu_4308_p2;
      sext_ln100_1_reg_4854 <= sext_ln100_1_fu_1596_p1;
      sext_ln100_reg_4849 <= sext_ln100_fu_1593_p1;
      sext_ln105_1_reg_4871 <= sext_ln105_1_fu_1599_p1;
      sext_ln111_1_reg_4896 <= sext_ln111_1_fu_1605_p1;
      sext_ln111_reg_4891 <= sext_ln111_fu_1602_p1;
      sext_ln91_reg_4810 <= sext_ln91_fu_1577_p1;
      sext_ln93_1_reg_4818 <= sext_ln93_1_fu_1584_p1;
      sext_ln96_1_reg_4836 <= sext_ln96_1_fu_1590_p1;
    end 
  end

  assign Const_185 = (1'd1 ^ working_key[442]);

  always @(posedge ap_clk) begin
    if(Const_185 == ap_CS_fsm_state22) begin
      mul_ln141_reg_5101 <= mul_ln141_fu_4509_p2;
      mul_ln142_reg_5106 <= mul_ln142_fu_4515_p2;
      sext_ln140_reg_5089 <= sext_ln140_fu_1882_p1;
    end 
  end

  assign Const_186 = (1'd0 ^ working_key[443]);
  assign Const_187 = (1'd1 ^ working_key[444]);
  assign Const_188 = (1'd0 ^ working_key[445]);

  always @(posedge ap_clk) begin
    if((Const_186 == ap_CS_fsm_state24) | (Const_187 == ap_CS_fsm_state22) | (Const_188 == ap_CS_fsm_state14)) begin
      reg_1114 <= L_ACF_q1;
      reg_1118 <= L_ACF_q0;
    end 
  end

  assign Const_189 = (1'd0 ^ working_key[446]);
  assign Const_190 = (1'd1 ^ working_key[447]);

  always @(posedge ap_clk) begin
    if((Const_189 == ap_CS_fsm_state48) | (Const_190 == ap_CS_fsm_state43)) begin
      reg_1122 <= P_q0;
    end 
  end

  assign Const_191 = (1'd0 ^ working_key[448]);
  assign Const_192 = (1'd0 ^ working_key[449]);
  assign Const_193 = (1'd0 ^ working_key[450]);

  always @(posedge ap_clk) begin
    if((Const_191 == and_ln72_reg_4687) & (icmp_ln75_fu_1524_p2 == Const_192) & (Const_193 == ap_CS_fsm_state6)) begin
      s_addr_2_reg_4709 <= zext_ln76_1_fu_1536_p1;
    end 
  end

  assign Const_194 = (1'd1 ^ working_key[451]);
  assign Const_195 = (1'd1 ^ working_key[452]);
  assign Const_196 = (1'd1 ^ working_key[453]);
  assign Const_197 = (1'd0 ^ working_key[454]);
  assign Const_198 = (1'd1 ^ working_key[455]);
  assign Const_199 = (1'd1 ^ working_key[456]);
  assign Const_200 = (1'd0 ^ working_key[457]);

  always @(posedge ap_clk) begin
    if((Const_194 == ap_CS_fsm_state44) & ((icmp_ln147_reg_5407 == Const_195) & (icmp_ln204_reg_5387 == Const_196) & (icmp_ln178_reg_5248 == Const_197) | (icmp_ln150_fu_2589_p2 == Const_198) & (icmp_ln204_reg_5387 == Const_199) & (icmp_ln178_reg_5248 == Const_200))) begin
      select_ln213_reg_5434 <= select_ln213_fu_2648_p3;
    end 
  end

  assign Const_201 = (1'd0 ^ working_key[458]);

  always @(posedge ap_clk) begin
    if(Const_201 == ap_CS_fsm_state52) begin
      select_ln273_reg_5552 <= select_ln273_fu_3151_p3;
    end 
  end

  assign Const_202 = (1'd1 ^ working_key[459]);

  always @(posedge ap_clk) begin
    if(Const_202 == ap_CS_fsm_state34) begin
      sext_ln187_reg_5292 <= sext_ln187_fu_2439_p1;
    end 
  end

  assign Const_203 = (1'd0 ^ working_key[460]);

  always @(posedge ap_clk) begin
    if(Const_203 == ap_CS_fsm_state11) begin
      sl_1_reg_4732 <= s_q0;
    end 
  end

  assign Const_204 = (1'd1 ^ working_key[461]);

  always @(posedge ap_clk) begin
    if(Const_204 == ap_CS_fsm_state12) begin
      sl_2_reg_4754 <= s_q0;
      sl_3_reg_4760 <= s_q1;
    end 
  end

  assign Const_205 = (1'd0 ^ working_key[462]);

  always @(posedge ap_clk) begin
    if(Const_205 == ap_CS_fsm_state13) begin
      sl_4_reg_4788 <= s_q1;
      sl_5_reg_4794 <= s_q0;
    end 
  end

  assign Const_206 = (1'd0 ^ working_key[463]);

  always @(posedge ap_clk) begin
    if(Const_206 == ap_CS_fsm_state46) begin
      sub_ln223_reg_5468 <= sub_ln223_fu_2782_p2;
    end 
  end

  assign Const_207 = (1'd1 ^ working_key[464]);

  always @(posedge ap_clk) begin
    if(Const_207 == ap_CS_fsm_state7) begin
      trunc_ln2_reg_4714 <= { { grp_fu_4288_p3[30:15] } };
    end 
  end

  assign Const_208 = (1'd1 ^ working_key[465]);
  assign Const_209 = (1'd0 ^ working_key[466]);

  always @(posedge ap_clk) begin
    if((Const_208 == and_ln72_fu_1495_p2) & (Const_209 == ap_CS_fsm_state4)) begin
      trunc_ln76_reg_4691 <= trunc_ln76_fu_1501_p1;
    end 
  end

  assign Const_210 = (1'd0 ^ working_key[467]);
  assign Const_211 = (1'd0 ^ working_key[468]);

  always @(posedge ap_clk) begin
    if((icmp_ln186_fu_2443_p2 == Const_210) & (Const_211 == ap_CS_fsm_state35)) begin
      zext_ln187_reg_5305[3:0] <= zext_ln187_fu_2455_p1[3:0];
    end 
  end

  assign Const_212 = (1'd1 ^ working_key[469]);
  assign Const_213 = (1'd0 ^ working_key[470]);

  always @(posedge ap_clk) begin
    if((icmp_ln194_fu_2497_p2 == Const_212) & (Const_213 == ap_CS_fsm_state39)) begin
      zext_ln195_reg_5341[3:0] <= zext_ln195_fu_2509_p1[3:0];
    end 
  end

  assign Const_214 = (1'd0 ^ working_key[471]);
  assign Const_215 = (1'd0 ^ working_key[472]);

  always @(posedge ap_clk) begin
    if((icmp_ln204_fu_2555_p2 == Const_214) & (Const_215 == ap_CS_fsm_state43)) begin
      zext_ln206_1_reg_5411[3:0] <= zext_ln206_1_fu_2579_p1[3:0];
    end 
  end

  assign Const_216 = (1'd0 ^ working_key[473]);

  always @(posedge ap_clk) begin
    if(Const_216 == ap_CS_fsm_state5) begin
      zext_ln75_reg_4696[14:0] <= zext_ln75_fu_1520_p1[14:0];
    end 
  end

  assign Const_217 = (1'd0 ^ working_key[474]);
  assign Const_218 = (1'd1 ^ working_key[475]);
  assign Const_219 = (1'd0 ^ working_key[476]);

  always @(*) begin
    if(((Const_217 == ap_CS_fsm_state39) ^ working_key[479]) == 1'b1) begin
      ACF_address0 = zext_ln195_fu_2509_p1;
    end else if(((Const_218 == ap_CS_fsm_state37) ^ working_key[478]) == 1'b0) begin
      ACF_address0 = zext_ln193_fu_2486_p1;
    end else if(((Const_219 == ap_CS_fsm_state36) ^ working_key[477]) == 1'b1) begin
      ACF_address0 = zext_ln187_reg_5305;
    end else begin
      ACF_address0 = 'bx;
    end
  end

  assign Const_220 = (1'd0 ^ working_key[480]);
  assign Const_221 = (1'd1 ^ working_key[481]);
  assign Const_222 = (1'd1 ^ working_key[482]);
  assign Const_223 = (1'd0 ^ working_key[483]);
  assign Const_224 = (1'd0 ^ working_key[484]);

  always @(*) begin
    if((((Const_220 == ap_CS_fsm_state36) | (Const_221 == ap_CS_fsm_state39) | (Const_222 == ap_CS_fsm_state37)) ^ working_key[485]) == 1'b1) begin
      ACF_ce0 = Const_224;
    end else begin
      ACF_ce0 = Const_223;
    end
  end

  assign Const_225 = (1'd1 ^ working_key[486]);
  assign Const_226 = (1'd0 ^ working_key[487]);
  assign Const_227 = (1'd0 ^ working_key[488]);

  always @(*) begin
    if(((Const_225 == ap_CS_fsm_state36) ^ working_key[489]) == 1'b1) begin
      ACF_we0 = Const_227;
    end else begin
      ACF_we0 = Const_226;
    end
  end

  assign Const_228 = (1'd1 ^ working_key[490]);
  assign Const_229 = (1'd0 ^ working_key[491]);
  assign Const_230 = (1'd1 ^ working_key[492]);

  always @(*) begin
    if(((Const_228 == ap_CS_fsm_state49) ^ working_key[495]) == 1'b0) begin
      K_address0 = K_addr_1_reg_5481;
    end else if(((Const_229 == ap_CS_fsm_state47) ^ working_key[494]) == 1'b1) begin
      K_address0 = zext_ln225_fu_2793_p1;
    end else if(((Const_230 == ap_CS_fsm_state38) ^ working_key[493]) == 1'b1) begin
      K_address0 = 'bx;
    end else begin
      K_address0 = zext_ln193_reg_5318;
    end
  end

  assign Const_231 = (1'd1 ^ working_key[496]);
  assign Const_232 = (1'd0 ^ working_key[497]);
  assign Const_233 = (1'd1 ^ working_key[498]);
  assign Const_234 = (1'd0 ^ working_key[499]);
  assign Const_235 = (1'd0 ^ working_key[500]);

  always @(*) begin
    if((((Const_231 == ap_CS_fsm_state49) | (Const_232 == ap_CS_fsm_state38) | (Const_233 == ap_CS_fsm_state47)) ^ working_key[501]) == 1'b1) begin
      K_ce0 = Const_235;
    end else begin
      K_ce0 = Const_234;
    end
  end

  assign Const_236 = (1'd1 ^ working_key[502]);
  assign Const_237 = (1'd1 ^ working_key[503]);

  always @(*) begin
    if(((Const_236 == ap_CS_fsm_state49) ^ working_key[505]) == 1'b1) begin
      K_d0 = select_ln40_5_fu_2994_p3;
    end else if(((Const_237 == ap_CS_fsm_state38) ^ working_key[504]) == 1'b1) begin
      K_d0 = ACF_q0;
    end else begin
      K_d0 = 'bx;
    end
  end

  assign Const_238 = (1'd1 ^ working_key[506]);
  assign Const_239 = (1'd0 ^ working_key[507]);
  assign Const_240 = (1'd1 ^ working_key[508]);
  assign Const_241 = (1'd1 ^ working_key[509]);

  always @(*) begin
    if((((Const_238 == ap_CS_fsm_state49) | (Const_239 == ap_CS_fsm_state38)) ^ working_key[510]) == 1'b1) begin
      K_we0 = Const_240;
    end else begin
      K_we0 = Const_241;
    end
  end

  assign Const_242 = (1'd0 ^ working_key[511]);
  assign Const_243 = (1'd1 ^ working_key[512]);
  assign Const_244 = (1'd0 ^ working_key[513]);
  assign Const_245 = (1'd1 ^ working_key[514]);
  assign Const_246 = (3'd4 ^ working_key[517:515]);
  assign Const_247 = (1'd1 ^ working_key[518]);
  assign Const_248 = (3'd2 ^ working_key[521:519]);
  assign Const_249 = (1'd1 ^ working_key[522]);
  assign Const_250 = (3'd0 ^ working_key[525:523]);
  assign Const_251 = (1'd1 ^ working_key[526]);
  assign Const_252 = (3'd2 ^ working_key[529:527]);
  assign Const_253 = (1'd0 ^ working_key[530]);
  assign Const_254 = (1'd0 ^ working_key[531]);
  assign Const_255 = (3'd6 ^ working_key[534:532]);
  assign Const_256 = (1'd1 ^ working_key[535]);
  assign Const_257 = (1'd0 ^ working_key[536]);
  assign Const_258 = (1'd0 ^ working_key[537]);
  assign Const_259 = (1'd0 ^ working_key[538]);
  assign Const_260 = (1'd1 ^ working_key[539]);
  assign Const_261 = (1'd1 ^ working_key[540]);
  assign Const_262 = (1'd1 ^ working_key[541]);
  assign Const_263 = (1'd0 ^ working_key[542]);
  assign Const_264 = (1'd1 ^ working_key[543]);
  assign Const_265 = (1'd1 ^ working_key[544]);
  assign Const_266 = (1'd1 ^ working_key[545]);
  assign Const_267 = (1'd1 ^ working_key[546]);
  assign Const_268 = (1'd1 ^ working_key[547]);
  assign Const_269 = (1'd0 ^ working_key[548]);

  always @(*) begin
    if(((Const_242 == ap_CS_fsm_state60) ^ working_key[560]) == 1'b1) begin
      LARc_address0 = LARc_addr_11_reg_5638;
    end else if(((Const_243 == ap_CS_fsm_state59) ^ working_key[559]) == 1'b0) begin
      LARc_address0 = LARc_addr_9_reg_5612;
    end else if(((Const_244 == ap_CS_fsm_state58) ^ working_key[558]) == 1'b1) begin
      LARc_address0 = LARc_addr_7_reg_5582;
    end else if(((Const_245 == ap_CS_fsm_state57) ^ working_key[557]) == 1'b0) begin
      LARc_address0 = Const_246;
    end else if(((Const_247 == ap_CS_fsm_state56) ^ working_key[556]) == 1'b1) begin
      LARc_address0 = Const_248;
    end else if(((Const_249 == ap_CS_fsm_state55) ^ working_key[555]) == 1'b0) begin
      LARc_address0 = Const_250;
    end else if(((Const_251 == ap_CS_fsm_state54) ^ working_key[554]) == 1'b1) begin
      LARc_address0 = Const_252;
    end else if(((icmp_ln253_fu_3025_p2 == Const_253) & (Const_254 == ap_CS_fsm_state51) ^ working_key[553]) == 1'b1) begin
      LARc_address0 = Const_255;
    end else if(((icmp_ln253_fu_3025_p2 == Const_256) & (Const_257 == ap_CS_fsm_state51) ^ working_key[552]) == 1'b0) begin
      LARc_address0 = p_0_rec_i16_cast_fu_3020_p1;
    end else if(((Const_258 == ap_CS_fsm_state50) ^ working_key[551]) == 1'b1) begin
      LARc_address0 = p_0_rec_i1_cast_fu_3003_p1;
    end else if(((icmp_ln204_reg_5387 == Const_259) & (icmp_ln206_fu_2677_p2 == Const_260) & (icmp_ln178_reg_5248 == Const_261) & (Const_262 == ap_CS_fsm_state44) ^ working_key[550]) == 1'b1) begin
      LARc_address0 = sum42_cast_fu_2672_p1;
    end else if(((Const_263 == ap_CS_fsm_state44) & ((icmp_ln147_reg_5407 == Const_264) & (icmp_ln204_reg_5387 == Const_265) & (icmp_ln178_reg_5248 == Const_266) | (icmp_ln150_fu_2589_p2 == Const_267) & (icmp_ln204_reg_5387 == Const_268) & (icmp_ln178_reg_5248 == Const_269)) ^ working_key[549]) == 1'b1) begin
      LARc_address0 = 'bx;
    end else begin
      LARc_address0 = LARc_addr_2_reg_5361;
    end
  end

  assign Const_270 = (1'd0 ^ working_key[561]);
  assign Const_271 = (1'd0 ^ working_key[562]);
  assign Const_272 = (1'd1 ^ working_key[563]);
  assign Const_273 = (1'd1 ^ working_key[564]);
  assign Const_274 = (3'd5 ^ working_key[567:565]);
  assign Const_275 = (1'd0 ^ working_key[568]);
  assign Const_276 = (3'd3 ^ working_key[571:569]);
  assign Const_277 = (1'd1 ^ working_key[572]);
  assign Const_278 = (3'd1 ^ working_key[575:573]);
  assign Const_279 = (1'd1 ^ working_key[576]);
  assign Const_280 = (3'd1 ^ working_key[579:577]);
  assign Const_281 = (1'd0 ^ working_key[580]);
  assign Const_282 = (1'd1 ^ working_key[581]);
  assign Const_283 = (3'd0 ^ working_key[584:582]);

  always @(*) begin
    if(((Const_270 == ap_CS_fsm_state60) ^ working_key[593]) == 1'b1) begin
      LARc_address1 = LARc_addr_10_reg_5633;
    end else if(((Const_271 == ap_CS_fsm_state59) ^ working_key[592]) == 1'b0) begin
      LARc_address1 = LARc_addr_8_reg_5607;
    end else if(((Const_272 == ap_CS_fsm_state58) ^ working_key[591]) == 1'b1) begin
      LARc_address1 = LARc_addr_6_reg_5577;
    end else if(((Const_273 == ap_CS_fsm_state57) ^ working_key[590]) == 1'b0) begin
      LARc_address1 = Const_274;
    end else if(((Const_275 == ap_CS_fsm_state56) ^ working_key[589]) == 1'b1) begin
      LARc_address1 = Const_276;
    end else if(((Const_277 == ap_CS_fsm_state55) ^ working_key[588]) == 1'b0) begin
      LARc_address1 = Const_278;
    end else if(((Const_279 == ap_CS_fsm_state54) ^ working_key[587]) == 1'b1) begin
      LARc_address1 = Const_280;
    end else if(((Const_281 == ap_CS_fsm_state53) ^ working_key[586]) == 1'b1) begin
      LARc_address1 = LARc_addr_4_reg_5532;
    end else if(((Const_282 == ap_CS_fsm_state51) ^ working_key[585]) == 1'b1) begin
      LARc_address1 = 'bx;
    end else begin
      LARc_address1 = Const_283;
    end
  end

  assign Const_284 = (1'd0 ^ working_key[594]);
  assign Const_285 = (1'd0 ^ working_key[595]);
  assign Const_286 = (1'd1 ^ working_key[596]);
  assign Const_287 = (1'd1 ^ working_key[597]);
  assign Const_288 = (1'd0 ^ working_key[598]);
  assign Const_289 = (1'd1 ^ working_key[599]);
  assign Const_290 = (1'd0 ^ working_key[600]);
  assign Const_291 = (1'd0 ^ working_key[601]);
  assign Const_292 = (1'd0 ^ working_key[602]);
  assign Const_293 = (1'd0 ^ working_key[603]);
  assign Const_294 = (1'd1 ^ working_key[604]);
  assign Const_295 = (1'd0 ^ working_key[605]);
  assign Const_296 = (1'd0 ^ working_key[606]);
  assign Const_297 = (1'd1 ^ working_key[607]);
  assign Const_298 = (1'd1 ^ working_key[608]);
  assign Const_299 = (1'd0 ^ working_key[609]);
  assign Const_300 = (1'd0 ^ working_key[610]);
  assign Const_301 = (1'd0 ^ working_key[611]);
  assign Const_302 = (1'd1 ^ working_key[612]);
  assign Const_303 = (1'd1 ^ working_key[613]);
  assign Const_304 = (1'd0 ^ working_key[614]);
  assign Const_305 = (1'd1 ^ working_key[615]);
  assign Const_306 = (1'd1 ^ working_key[616]);
  assign Const_307 = (1'd0 ^ working_key[617]);
  assign Const_308 = (1'd0 ^ working_key[618]);

  always @(*) begin
    if((((Const_284 == ap_CS_fsm_state58) | (Const_285 == ap_CS_fsm_state57) | (Const_286 == ap_CS_fsm_state56) | (Const_287 == ap_CS_fsm_state55) | (Const_288 == ap_CS_fsm_state54) | (Const_289 == ap_CS_fsm_state50) | (Const_290 == ap_CS_fsm_state60) | (Const_291 == ap_CS_fsm_state59) | (icmp_ln253_fu_3025_p2 == Const_292) & (Const_293 == ap_CS_fsm_state51) | (icmp_ln253_fu_3025_p2 == Const_294) & (Const_295 == ap_CS_fsm_state51) | (Const_296 == ap_CS_fsm_state44) & ((icmp_ln147_reg_5407 == Const_297) & (icmp_ln204_reg_5387 == Const_298) & (icmp_ln178_reg_5248 == Const_299) | (icmp_ln150_fu_2589_p2 == Const_300) & (icmp_ln204_reg_5387 == Const_301) & (icmp_ln178_reg_5248 == Const_302)) | (icmp_ln204_reg_5387 == Const_303) & (icmp_ln206_fu_2677_p2 == Const_304) & (icmp_ln178_reg_5248 == Const_305) & (Const_306 == ap_CS_fsm_state44)) ^ working_key[619]) == 1'b1) begin
      LARc_ce0 = Const_308;
    end else begin
      LARc_ce0 = Const_307;
    end
  end

  assign Const_309 = (1'd1 ^ working_key[620]);
  assign Const_310 = (1'd0 ^ working_key[621]);
  assign Const_311 = (1'd1 ^ working_key[622]);
  assign Const_312 = (1'd0 ^ working_key[623]);
  assign Const_313 = (1'd1 ^ working_key[624]);
  assign Const_314 = (1'd0 ^ working_key[625]);
  assign Const_315 = (1'd1 ^ working_key[626]);
  assign Const_316 = (1'd0 ^ working_key[627]);
  assign Const_317 = (1'd1 ^ working_key[628]);
  assign Const_318 = (1'd0 ^ working_key[629]);
  assign Const_319 = (1'd0 ^ working_key[630]);

  always @(*) begin
    if((((Const_309 == ap_CS_fsm_state53) | (Const_310 == ap_CS_fsm_state58) | (Const_311 == ap_CS_fsm_state57) | (Const_312 == ap_CS_fsm_state56) | (Const_313 == ap_CS_fsm_state55) | (Const_314 == ap_CS_fsm_state54) | (Const_315 == ap_CS_fsm_state51) | (Const_316 == ap_CS_fsm_state60) | (Const_317 == ap_CS_fsm_state59)) ^ working_key[631]) == 1'b1) begin
      LARc_ce1 = Const_319;
    end else begin
      LARc_ce1 = Const_318;
    end
  end

  assign Const_320 = (1'd1 ^ working_key[632]);
  assign Const_321 = (1'd0 ^ working_key[633]);
  assign Const_322 = (1'd1 ^ working_key[634]);
  assign Const_323 = (1'd1 ^ working_key[635]);
  assign Const_324 = (1'd1 ^ working_key[636]);
  assign Const_325 = (1'd1 ^ working_key[637]);
  assign Const_326 = (1'd0 ^ working_key[638]);
  assign Const_327 = (1'd1 ^ working_key[639]);
  assign Const_328 = (1'd1 ^ working_key[640]);
  assign Const_329 = (16'd21845 ^ working_key[656:641]);
  assign Const_330 = (1'd0 ^ working_key[657]);
  assign Const_331 = (1'd1 ^ working_key[658]);
  assign Const_332 = (1'd1 ^ working_key[659]);
  assign Const_333 = (1'd0 ^ working_key[660]);
  assign Const_334 = (1'd1 ^ working_key[661]);
  assign Const_335 = (1'd1 ^ working_key[662]);
  assign Const_336 = (1'd1 ^ working_key[663]);

  always @(*) begin
    if(((Const_320 == ap_CS_fsm_state60) ^ working_key[669]) == 1'b1) begin
      LARc_d0 = sext_ln312_1_fu_4283_p1;
    end else if(((Const_321 == ap_CS_fsm_state59) ^ working_key[668]) == 1'b0) begin
      LARc_d0 = sext_ln310_1_fu_4153_p1;
    end else if(((Const_322 == ap_CS_fsm_state58) ^ working_key[667]) == 1'b1) begin
      LARc_d0 = sext_ln307_1_fu_3963_p1;
    end else if(((Const_323 == ap_CS_fsm_state57) ^ working_key[666]) == 1'b0) begin
      LARc_d0 = sext_ln305_1_fu_3727_p1;
    end else if((((Const_324 == ap_CS_fsm_state50) | (icmp_ln204_reg_5387 == Const_325) & (icmp_ln206_fu_2677_p2 == Const_326) & (icmp_ln178_reg_5248 == Const_327) & (Const_328 == ap_CS_fsm_state44)) ^ working_key[665]) == 1'b1) begin
      LARc_d0 = Const_329;
    end else if(((Const_330 == ap_CS_fsm_state44) & ((icmp_ln147_reg_5407 == Const_331) & (icmp_ln204_reg_5387 == Const_332) & (icmp_ln178_reg_5248 == Const_333) | (icmp_ln150_fu_2589_p2 == Const_334) & (icmp_ln204_reg_5387 == Const_335) & (icmp_ln178_reg_5248 == Const_336)) ^ working_key[664]) == 1'b1) begin
      LARc_d0 = select_ln213_fu_2648_p3;
    end else begin
      LARc_d0 = 'bx;
    end
  end

  assign Const_337 = (1'd0 ^ working_key[670]);
  assign Const_338 = (1'd1 ^ working_key[671]);
  assign Const_339 = (1'd0 ^ working_key[672]);
  assign Const_340 = (1'd0 ^ working_key[673]);
  assign Const_341 = (1'd1 ^ working_key[674]);

  always @(*) begin
    if(((Const_337 == ap_CS_fsm_state60) ^ working_key[679]) == 1'b1) begin
      LARc_d1 = sext_ln311_1_fu_4218_p1;
    end else if(((Const_338 == ap_CS_fsm_state59) ^ working_key[678]) == 1'b1) begin
      LARc_d1 = sext_ln309_1_fu_4088_p1;
    end else if(((Const_339 == ap_CS_fsm_state58) ^ working_key[677]) == 1'b0) begin
      LARc_d1 = sext_ln306_1_fu_3898_p1;
    end else if(((Const_340 == ap_CS_fsm_state57) ^ working_key[676]) == 1'b1) begin
      LARc_d1 = sext_ln304_1_fu_3662_p1;
    end else if(((Const_341 == ap_CS_fsm_state53) ^ working_key[675]) == 1'b1) begin
      LARc_d1 = 'bx;
    end else begin
      LARc_d1 = select_ln273_reg_5552;
    end
  end

  assign Const_342 = (1'd0 ^ working_key[680]);
  assign Const_343 = (1'd1 ^ working_key[681]);
  assign Const_344 = (1'd1 ^ working_key[682]);
  assign Const_345 = (1'd0 ^ working_key[683]);
  assign Const_346 = (1'd0 ^ working_key[684]);
  assign Const_347 = (1'd0 ^ working_key[685]);
  assign Const_348 = (1'd1 ^ working_key[686]);
  assign Const_349 = (1'd0 ^ working_key[687]);
  assign Const_350 = (1'd0 ^ working_key[688]);
  assign Const_351 = (1'd1 ^ working_key[689]);
  assign Const_352 = (1'd0 ^ working_key[690]);
  assign Const_353 = (1'd0 ^ working_key[691]);
  assign Const_354 = (1'd0 ^ working_key[692]);
  assign Const_355 = (1'd0 ^ working_key[693]);
  assign Const_356 = (1'd0 ^ working_key[694]);
  assign Const_357 = (1'd1 ^ working_key[695]);
  assign Const_358 = (1'd0 ^ working_key[696]);
  assign Const_359 = (1'd0 ^ working_key[697]);
  assign Const_360 = (1'd0 ^ working_key[698]);

  always @(*) begin
    if((((Const_342 == ap_CS_fsm_state58) | (Const_343 == ap_CS_fsm_state57) | (Const_344 == ap_CS_fsm_state60) | (Const_345 == ap_CS_fsm_state59) | (icmp_ln180_fu_3008_p2 == Const_346) & (Const_347 == ap_CS_fsm_state50) | (Const_348 == ap_CS_fsm_state44) & ((icmp_ln147_reg_5407 == Const_349) & (icmp_ln204_reg_5387 == Const_350) & (icmp_ln178_reg_5248 == Const_351) | (icmp_ln150_fu_2589_p2 == Const_352) & (icmp_ln204_reg_5387 == Const_353) & (icmp_ln178_reg_5248 == Const_354)) | (icmp_ln204_reg_5387 == Const_355) & (icmp_ln206_fu_2677_p2 == Const_356) & (icmp_ln178_reg_5248 == Const_357) & (Const_358 == ap_CS_fsm_state44)) ^ working_key[699]) == 1'b1) begin
      LARc_we0 = Const_360;
    end else begin
      LARc_we0 = Const_359;
    end
  end

  assign Const_361 = (1'd1 ^ working_key[700]);
  assign Const_362 = (1'd0 ^ working_key[701]);
  assign Const_363 = (1'd1 ^ working_key[702]);
  assign Const_364 = (1'd0 ^ working_key[703]);
  assign Const_365 = (1'd1 ^ working_key[704]);
  assign Const_366 = (1'd0 ^ working_key[705]);
  assign Const_367 = (1'd1 ^ working_key[706]);

  always @(*) begin
    if((((Const_361 == ap_CS_fsm_state53) | (Const_362 == ap_CS_fsm_state58) | (Const_363 == ap_CS_fsm_state57) | (Const_364 == ap_CS_fsm_state60) | (Const_365 == ap_CS_fsm_state59)) ^ working_key[707]) == 1'b1) begin
      LARc_we1 = Const_366;
    end else begin
      LARc_we1 = Const_367;
    end
  end

  assign Const_368 = (1'd0 ^ working_key[708]);
  assign Const_369 = (1'd1 ^ working_key[709]);
  assign Const_370 = (4'd1 ^ working_key[713:710]);
  assign Const_371 = (1'd1 ^ working_key[714]);
  assign Const_372 = (4'd12 ^ working_key[718:715]);
  assign Const_373 = (1'd1 ^ working_key[719]);
  assign Const_374 = (4'd9 ^ working_key[723:720]);
  assign Const_375 = (1'd1 ^ working_key[724]);
  assign Const_376 = (4'd8 ^ working_key[728:725]);
  assign Const_377 = (1'd0 ^ working_key[729]);
  assign Const_378 = (1'd0 ^ working_key[730]);
  assign Const_379 = (1'd0 ^ working_key[731]);
  assign Const_380 = (1'd0 ^ working_key[732]);
  assign Const_381 = (1'd0 ^ working_key[733]);
  assign Const_382 = (1'd0 ^ working_key[734]);
  assign Const_383 = (1'd1 ^ working_key[735]);
  assign Const_384 = (1'd0 ^ working_key[736]);
  assign Const_385 = (4'd11 ^ working_key[740:737]);
  assign Const_386 = (1'd1 ^ working_key[741]);
  assign Const_387 = (4'd13 ^ working_key[745:742]);
  assign Const_388 = (1'd1 ^ working_key[746]);
  assign Const_389 = (4'd0 ^ working_key[750:747]);
  assign Const_390 = (1'd0 ^ working_key[751]);
  assign Const_391 = (4'd9 ^ working_key[755:752]);
  assign Const_392 = (1'd1 ^ working_key[756]);
  assign Const_393 = (1'd0 ^ working_key[757]);
  assign Const_394 = (4'd10 ^ working_key[761:758]);
  assign Const_395 = (1'd1 ^ working_key[762]);

  always @(*) begin
    if(((Const_368 == ap_CS_fsm_state29) ^ working_key[776]) == 1'b1) begin
      L_ACF_address0 = zext_ln152_fu_2060_p1;
    end else if(((Const_369 == ap_CS_fsm_state23) ^ working_key[775]) == 1'b0) begin
      L_ACF_address0 = Const_370;
    end else if(((Const_371 == ap_CS_fsm_state22) ^ working_key[774]) == 1'b1) begin
      L_ACF_address0 = Const_372;
    end else if(((Const_373 == ap_CS_fsm_state21) ^ working_key[773]) == 1'b0) begin
      L_ACF_address0 = Const_374;
    end else if(((Const_375 == ap_CS_fsm_state20) ^ working_key[772]) == 1'b1) begin
      L_ACF_address0 = Const_376;
    end else if((((Const_377 == ap_CS_fsm_state19) | (Const_378 == ap_CS_fsm_state27)) ^ working_key[771]) == 1'b0) begin
      L_ACF_address0 = L_ACF_addr_7_reg_5023;
    end else if((((Const_379 == ap_CS_fsm_state26) | (Const_380 == ap_CS_fsm_state18)) ^ working_key[770]) == 1'b1) begin
      L_ACF_address0 = L_ACF_addr_5_reg_4911;
    end else if((((Const_381 == ap_CS_fsm_state25) | (Const_382 == ap_CS_fsm_state17)) ^ working_key[769]) == 1'b0) begin
      L_ACF_address0 = L_ACF_addr_3_reg_4782;
    end else if((((Const_383 == ap_CS_fsm_state16) | (Const_384 == ap_CS_fsm_state24)) ^ working_key[768]) == 1'b1) begin
      L_ACF_address0 = Const_385;
    end else if(((Const_386 == ap_CS_fsm_state15) ^ working_key[767]) == 1'b0) begin
      L_ACF_address0 = Const_387;
    end else if(((Const_388 == ap_CS_fsm_state14) ^ working_key[766]) == 1'b1) begin
      L_ACF_address0 = Const_389;
    end else if(((Const_390 == ap_CS_fsm_state13) ^ working_key[765]) == 1'b1) begin
      L_ACF_address0 = Const_391;
    end else if((((Const_392 == ap_CS_fsm_state31) | (Const_393 == ap_CS_fsm_state12)) ^ working_key[764]) == 1'b1) begin
      L_ACF_address0 = Const_394;
    end else if(((Const_395 == ap_CS_fsm_state10) ^ working_key[763]) == 1'b1) begin
      L_ACF_address0 = zext_ln89_fu_1566_p1;
    end else begin
      L_ACF_address0 = 'bx;
    end
  end

  assign Const_396 = (1'd0 ^ working_key[777]);
  assign Const_397 = (1'd1 ^ working_key[778]);
  assign Const_398 = (1'd0 ^ working_key[779]);
  assign Const_399 = (4'd2 ^ working_key[783:780]);
  assign Const_400 = (1'd1 ^ working_key[784]);
  assign Const_401 = (4'd2 ^ working_key[788:785]);
  assign Const_402 = (1'd1 ^ working_key[789]);
  assign Const_403 = (4'd14 ^ working_key[793:790]);
  assign Const_404 = (1'd0 ^ working_key[794]);
  assign Const_405 = (4'd8 ^ working_key[798:795]);
  assign Const_406 = (1'd1 ^ working_key[799]);
  assign Const_407 = (1'd0 ^ working_key[800]);
  assign Const_408 = (1'd0 ^ working_key[801]);
  assign Const_409 = (1'd1 ^ working_key[802]);
  assign Const_410 = (1'd0 ^ working_key[803]);
  assign Const_411 = (1'd1 ^ working_key[804]);
  assign Const_412 = (1'd0 ^ working_key[805]);
  assign Const_413 = (1'd1 ^ working_key[806]);
  assign Const_414 = (1'd1 ^ working_key[807]);
  assign Const_415 = (4'd9 ^ working_key[811:808]);
  assign Const_416 = (1'd1 ^ working_key[812]);
  assign Const_417 = (4'd3 ^ working_key[816:813]);
  assign Const_418 = (1'd0 ^ working_key[817]);
  assign Const_419 = (4'd13 ^ working_key[821:818]);
  assign Const_420 = (1'd1 ^ working_key[822]);
  assign Const_421 = (4'd5 ^ working_key[826:823]);
  assign Const_422 = (1'd0 ^ working_key[827]);
  assign Const_423 = (4'd11 ^ working_key[831:828]);

  always @(*) begin
    if(((Const_396 == ap_CS_fsm_state35) ^ working_key[846]) == 1'b0) begin
      L_ACF_address1 = zext_ln187_fu_2455_p1;
    end else if(((Const_397 == ap_CS_fsm_state30) ^ working_key[845]) == 1'b1) begin
      L_ACF_address1 = L_ACF_addr_9_reg_5224;
    end else if(((Const_398 == ap_CS_fsm_state28) ^ working_key[844]) == 1'b0) begin
      L_ACF_address1 = Const_399;
    end else if(((Const_400 == ap_CS_fsm_state23) ^ working_key[843]) == 1'b1) begin
      L_ACF_address1 = Const_401;
    end else if(((Const_402 == ap_CS_fsm_state22) ^ working_key[842]) == 1'b1) begin
      L_ACF_address1 = Const_403;
    end else if(((Const_404 == ap_CS_fsm_state21) ^ working_key[841]) == 1'b0) begin
      L_ACF_address1 = Const_405;
    end else if(((Const_406 == ap_CS_fsm_state20) ^ working_key[840]) == 1'b1) begin
      L_ACF_address1 = L_ACF_addr_1_reg_4748;
    end else if((((Const_407 == ap_CS_fsm_state19) | (Const_408 == ap_CS_fsm_state27)) ^ working_key[839]) == 1'b1) begin
      L_ACF_address1 = L_ACF_addr_6_reg_4967;
    end else if((((Const_409 == ap_CS_fsm_state26) | (Const_410 == ap_CS_fsm_state18)) ^ working_key[838]) == 1'b0) begin
      L_ACF_address1 = L_ACF_addr_4_reg_4885;
    end else if((((Const_411 == ap_CS_fsm_state25) | (Const_412 == ap_CS_fsm_state17)) ^ working_key[837]) == 1'b1) begin
      L_ACF_address1 = L_ACF_addr_2_reg_4776;
    end else if((((Const_413 == ap_CS_fsm_state16) | (Const_414 == ap_CS_fsm_state24)) ^ working_key[836]) == 1'b0) begin
      L_ACF_address1 = Const_415;
    end else if(((Const_416 == ap_CS_fsm_state15) ^ working_key[835]) == 1'b1) begin
      L_ACF_address1 = Const_417;
    end else if(((Const_418 == ap_CS_fsm_state14) ^ working_key[834]) == 1'b0) begin
      L_ACF_address1 = Const_419;
    end else if(((Const_420 == ap_CS_fsm_state13) ^ working_key[833]) == 1'b0) begin
      L_ACF_address1 = Const_421;
    end else if(((Const_422 == ap_CS_fsm_state12) ^ working_key[832]) == 1'b1) begin
      L_ACF_address1 = Const_423;
    end else begin
      L_ACF_address1 = 'bx;
    end
  end

  assign Const_424 = (1'd1 ^ working_key[847]);
  assign Const_425 = (1'd0 ^ working_key[848]);
  assign Const_426 = (1'd1 ^ working_key[849]);
  assign Const_427 = (1'd0 ^ working_key[850]);
  assign Const_428 = (1'd0 ^ working_key[851]);
  assign Const_429 = (1'd1 ^ working_key[852]);
  assign Const_430 = (1'd1 ^ working_key[853]);
  assign Const_431 = (1'd0 ^ working_key[854]);
  assign Const_432 = (1'd1 ^ working_key[855]);
  assign Const_433 = (1'd0 ^ working_key[856]);
  assign Const_434 = (1'd0 ^ working_key[857]);
  assign Const_435 = (1'd0 ^ working_key[858]);
  assign Const_436 = (1'd0 ^ working_key[859]);
  assign Const_437 = (1'd0 ^ working_key[860]);
  assign Const_438 = (1'd0 ^ working_key[861]);
  assign Const_439 = (1'd0 ^ working_key[862]);
  assign Const_440 = (1'd1 ^ working_key[863]);
  assign Const_441 = (1'd0 ^ working_key[864]);
  assign Const_442 = (1'd1 ^ working_key[865]);
  assign Const_443 = (1'd0 ^ working_key[866]);
  assign Const_444 = (1'd0 ^ working_key[867]);

  always @(*) begin
    if((((Const_424 == ap_CS_fsm_state31) | (Const_425 == ap_CS_fsm_state29) | (Const_426 == ap_CS_fsm_state26) | (Const_427 == ap_CS_fsm_state25) | (Const_428 == ap_CS_fsm_state20) | (Const_429 == ap_CS_fsm_state19) | (Const_430 == ap_CS_fsm_state16) | (Const_431 == ap_CS_fsm_state12) | (Const_432 == ap_CS_fsm_state10) | (Const_433 == ap_CS_fsm_state24) | (Const_434 == ap_CS_fsm_state22) | (Const_435 == ap_CS_fsm_state15) | (Const_436 == ap_CS_fsm_state23) | (Const_437 == ap_CS_fsm_state13) | (Const_438 == ap_CS_fsm_state21) | (Const_439 == ap_CS_fsm_state14) | (Const_440 == ap_CS_fsm_state27) | (Const_441 == ap_CS_fsm_state18) | (Const_442 == ap_CS_fsm_state17)) ^ working_key[868]) == 1'b1) begin
      L_ACF_ce0 = Const_444;
    end else begin
      L_ACF_ce0 = Const_443;
    end
  end

  assign Const_445 = (1'd1 ^ working_key[869]);
  assign Const_446 = (1'd1 ^ working_key[870]);
  assign Const_447 = (1'd0 ^ working_key[871]);
  assign Const_448 = (1'd1 ^ working_key[872]);
  assign Const_449 = (1'd0 ^ working_key[873]);
  assign Const_450 = (1'd1 ^ working_key[874]);
  assign Const_451 = (1'd0 ^ working_key[875]);
  assign Const_452 = (1'd1 ^ working_key[876]);
  assign Const_453 = (1'd0 ^ working_key[877]);
  assign Const_454 = (1'd1 ^ working_key[878]);
  assign Const_455 = (1'd0 ^ working_key[879]);
  assign Const_456 = (1'd1 ^ working_key[880]);
  assign Const_457 = (1'd0 ^ working_key[881]);
  assign Const_458 = (1'd1 ^ working_key[882]);
  assign Const_459 = (1'd0 ^ working_key[883]);
  assign Const_460 = (1'd1 ^ working_key[884]);
  assign Const_461 = (1'd0 ^ working_key[885]);
  assign Const_462 = (1'd1 ^ working_key[886]);
  assign Const_463 = (1'd0 ^ working_key[887]);
  assign Const_464 = (1'd1 ^ working_key[888]);
  assign Const_465 = (1'd1 ^ working_key[889]);

  always @(*) begin
    if((((Const_445 == ap_CS_fsm_state30) | (Const_446 == ap_CS_fsm_state28) | (Const_447 == ap_CS_fsm_state35) | (Const_448 == ap_CS_fsm_state26) | (Const_449 == ap_CS_fsm_state25) | (Const_450 == ap_CS_fsm_state20) | (Const_451 == ap_CS_fsm_state19) | (Const_452 == ap_CS_fsm_state16) | (Const_453 == ap_CS_fsm_state12) | (Const_454 == ap_CS_fsm_state24) | (Const_455 == ap_CS_fsm_state22) | (Const_456 == ap_CS_fsm_state15) | (Const_457 == ap_CS_fsm_state23) | (Const_458 == ap_CS_fsm_state13) | (Const_459 == ap_CS_fsm_state21) | (Const_460 == ap_CS_fsm_state14) | (Const_461 == ap_CS_fsm_state27) | (Const_462 == ap_CS_fsm_state18) | (Const_463 == ap_CS_fsm_state17)) ^ working_key[890]) == 1'b1) begin
      L_ACF_ce1 = Const_464;
    end else begin
      L_ACF_ce1 = Const_465;
    end
  end

  assign Const_466 = (1'd1 ^ working_key[891]);
  assign Const_467 = (1'd1 ^ working_key[892]);
  assign Const_468 = (1'd1 ^ working_key[893]);
  assign Const_469 = (1'd1 ^ working_key[894]);
  assign Const_470 = (1'd0 ^ working_key[895]);
  assign Const_471 = (1'd1 ^ working_key[896]);
  assign Const_472 = (1'd0 ^ working_key[897]);
  assign Const_473 = (1'd1 ^ working_key[898]);
  assign Const_474 = (1'd0 ^ working_key[899]);
  assign Const_475 = (64'd7690576492028013226 ^ working_key[963:900]);

  always @(*) begin
    if(((Const_466 == ap_CS_fsm_state27) ^ working_key[972]) == 1'b0) begin
      L_ACF_d0 = add_ln147_reg_5211;
    end else if(((Const_467 == ap_CS_fsm_state26) ^ working_key[971]) == 1'b1) begin
      L_ACF_d0 = add_ln145_1_reg_5191;
    end else if(((Const_468 == ap_CS_fsm_state25) ^ working_key[970]) == 1'b1) begin
      L_ACF_d0 = add_ln143_1_reg_5161;
    end else if(((Const_469 == ap_CS_fsm_state24) ^ working_key[969]) == 1'b0) begin
      L_ACF_d0 = add_ln141_reg_5126;
    end else if(((Const_470 == ap_CS_fsm_state19) ^ working_key[968]) == 1'b1) begin
      L_ACF_d0 = add_ln133_reg_5049;
    end else if(((Const_471 == ap_CS_fsm_state18) ^ working_key[967]) == 1'b1) begin
      L_ACF_d0 = add_ln131_reg_5008;
    end else if(((Const_472 == ap_CS_fsm_state17) ^ working_key[966]) == 1'b0) begin
      L_ACF_d0 = add_ln129_reg_5034;
    end else if(((Const_473 == ap_CS_fsm_state16) ^ working_key[965]) == 1'b1) begin
      L_ACF_d0 = add_ln127_reg_4983;
    end else if(((Const_474 == ap_CS_fsm_state10) ^ working_key[964]) == 1'b1) begin
      L_ACF_d0 = 'bx;
    end else begin
      L_ACF_d0 = Const_475;
    end
  end

  assign Const_476 = (1'd1 ^ working_key[973]);
  assign Const_477 = (1'd0 ^ working_key[974]);
  assign Const_478 = (1'd1 ^ working_key[975]);
  assign Const_479 = (1'd0 ^ working_key[976]);
  assign Const_480 = (1'd1 ^ working_key[977]);
  assign Const_481 = (1'd0 ^ working_key[978]);
  assign Const_482 = (1'd0 ^ working_key[979]);
  assign Const_483 = (1'd1 ^ working_key[980]);
  assign Const_484 = (1'd1 ^ working_key[981]);
  assign Const_485 = (1'd0 ^ working_key[982]);

  always @(*) begin
    if(((Const_476 == ap_CS_fsm_state30) ^ working_key[992]) == 1'b0) begin
      L_ACF_d1 = shl_ln152_fu_2071_p2;
    end else if(((Const_477 == ap_CS_fsm_state28) ^ working_key[991]) == 1'b1) begin
      L_ACF_d1 = add_ln148_reg_5216;
    end else if(((Const_478 == ap_CS_fsm_state27) ^ working_key[990]) == 1'b0) begin
      L_ACF_d1 = add_ln146_1_reg_5196;
    end else if(((Const_479 == ap_CS_fsm_state26) ^ working_key[989]) == 1'b0) begin
      L_ACF_d1 = add_ln144_1_reg_5166;
    end else if(((Const_480 == ap_CS_fsm_state25) ^ working_key[988]) == 1'b0) begin
      L_ACF_d1 = add_ln142_1_reg_5131;
    end else if(((Const_481 == ap_CS_fsm_state24) ^ working_key[987]) == 1'b0) begin
      L_ACF_d1 = add_ln140_fu_1971_p2;
    end else if(((Const_482 == ap_CS_fsm_state19) ^ working_key[986]) == 1'b0) begin
      L_ACF_d1 = add_ln132_reg_5044;
    end else if(((Const_483 == ap_CS_fsm_state18) ^ working_key[985]) == 1'b0) begin
      L_ACF_d1 = add_ln130_reg_5039;
    end else if(((Const_484 == ap_CS_fsm_state17) ^ working_key[984]) == 1'b0) begin
      L_ACF_d1 = add_ln128_reg_4988;
    end else if(((Const_485 == ap_CS_fsm_state16) ^ working_key[983]) == 1'b1) begin
      L_ACF_d1 = add_ln126_fu_1775_p2;
    end else begin
      L_ACF_d1 = 'bx;
    end
  end

  assign Const_486 = (1'd1 ^ working_key[993]);
  assign Const_487 = (1'd0 ^ working_key[994]);
  assign Const_488 = (1'd1 ^ working_key[995]);
  assign Const_489 = (1'd0 ^ working_key[996]);
  assign Const_490 = (1'd1 ^ working_key[997]);
  assign Const_491 = (1'd1 ^ working_key[998]);
  assign Const_492 = (1'd0 ^ working_key[999]);
  assign Const_493 = (1'd1 ^ working_key[1000]);
  assign Const_494 = (1'd1 ^ working_key[1001]);
  assign Const_495 = (1'd1 ^ working_key[1002]);
  assign Const_496 = (1'd0 ^ working_key[1003]);
  assign Const_497 = (1'd0 ^ working_key[1004]);

  always @(*) begin
    if((((Const_486 == ap_CS_fsm_state26) | (Const_487 == ap_CS_fsm_state25) | (Const_488 == ap_CS_fsm_state19) | (Const_489 == ap_CS_fsm_state16) | (Const_490 == ap_CS_fsm_state24) | (Const_491 == ap_CS_fsm_state27) | (Const_492 == ap_CS_fsm_state18) | (Const_493 == ap_CS_fsm_state17) | (tmp_14_fu_1558_p3 == Const_494) & (Const_495 == ap_CS_fsm_state10)) ^ working_key[1005]) == 1'b1) begin
      L_ACF_we0 = Const_497;
    end else begin
      L_ACF_we0 = Const_496;
    end
  end

  assign Const_498 = (1'd1 ^ working_key[1006]);
  assign Const_499 = (1'd0 ^ working_key[1007]);
  assign Const_500 = (1'd1 ^ working_key[1008]);
  assign Const_501 = (1'd0 ^ working_key[1009]);
  assign Const_502 = (1'd1 ^ working_key[1010]);
  assign Const_503 = (1'd0 ^ working_key[1011]);
  assign Const_504 = (1'd1 ^ working_key[1012]);
  assign Const_505 = (1'd0 ^ working_key[1013]);
  assign Const_506 = (1'd1 ^ working_key[1014]);
  assign Const_507 = (1'd0 ^ working_key[1015]);
  assign Const_508 = (1'd1 ^ working_key[1016]);
  assign Const_509 = (1'd1 ^ working_key[1017]);

  always @(*) begin
    if((((Const_498 == ap_CS_fsm_state30) | (Const_499 == ap_CS_fsm_state28) | (Const_500 == ap_CS_fsm_state26) | (Const_501 == ap_CS_fsm_state25) | (Const_502 == ap_CS_fsm_state19) | (Const_503 == ap_CS_fsm_state16) | (Const_504 == ap_CS_fsm_state24) | (Const_505 == ap_CS_fsm_state27) | (Const_506 == ap_CS_fsm_state18) | (Const_507 == ap_CS_fsm_state17)) ^ working_key[1018]) == 1'b1) begin
      L_ACF_we1 = Const_508;
    end else begin
      L_ACF_we1 = Const_509;
    end
  end

  assign Const_510 = (1'd1 ^ working_key[1019]);
  assign Const_511 = (1'd1 ^ working_key[1020]);
  assign Const_512 = (1'd1 ^ working_key[1021]);
  assign Const_513 = (1'd1 ^ working_key[1022]);
  assign Const_514 = (4'd5 ^ working_key[1026:1023]);
  assign Const_515 = (1'd0 ^ working_key[1027]);
  assign Const_516 = (4'd11 ^ working_key[1031:1028]);
  assign Const_517 = (1'd1 ^ working_key[1032]);

  always @(*) begin
    if(((Const_510 == ap_CS_fsm_state49) ^ working_key[1037]) == 1'b0) begin
      P_address0 = zext_ln225_reg_5476;
    end else if(((Const_511 == ap_CS_fsm_state47) ^ working_key[1036]) == 1'b1) begin
      P_address0 = zext_ln226_fu_2804_p1;
    end else if((((Const_512 == ap_CS_fsm_state46) | (Const_513 == ap_CS_fsm_state42)) ^ working_key[1035]) == 1'b0) begin
      P_address0 = Const_514;
    end else if(((Const_515 == ap_CS_fsm_state41) ^ working_key[1034]) == 1'b1) begin
      P_address0 = Const_516;
    end else if(((Const_517 == ap_CS_fsm_state40) ^ working_key[1033]) == 1'b1) begin
      P_address0 = 'bx;
    end else begin
      P_address0 = zext_ln195_reg_5341;
    end
  end

  assign Const_518 = (1'd1 ^ working_key[1038]);
  assign Const_519 = (1'd0 ^ working_key[1039]);
  assign Const_520 = (1'd1 ^ working_key[1040]);
  assign Const_521 = (1'd0 ^ working_key[1041]);
  assign Const_522 = (1'd1 ^ working_key[1042]);
  assign Const_523 = (1'd0 ^ working_key[1043]);
  assign Const_524 = (1'd1 ^ working_key[1044]);
  assign Const_525 = (1'd0 ^ working_key[1045]);

  always @(*) begin
    if((((Const_518 == ap_CS_fsm_state49) | (Const_519 == ap_CS_fsm_state40) | (Const_520 == ap_CS_fsm_state47) | (Const_521 == ap_CS_fsm_state46) | (Const_522 == ap_CS_fsm_state42) | (Const_523 == ap_CS_fsm_state41)) ^ working_key[1046]) == 1'b1) begin
      P_ce0 = Const_525;
    end else begin
      P_ce0 = Const_524;
    end
  end

  assign Const_526 = (1'd0 ^ working_key[1047]);
  assign Const_527 = (1'd1 ^ working_key[1048]);
  assign Const_528 = (1'd1 ^ working_key[1049]);

  always @(*) begin
    if(((Const_526 == ap_CS_fsm_state49) ^ working_key[1052]) == 1'b0) begin
      P_d0 = select_ln40_3_fu_2936_p3;
    end else if(((Const_527 == ap_CS_fsm_state46) ^ working_key[1051]) == 1'b1) begin
      P_d0 = select_ln40_1_reg_5463;
    end else if(((Const_528 == ap_CS_fsm_state40) ^ working_key[1050]) == 1'b1) begin
      P_d0 = 'bx;
    end else begin
      P_d0 = ACF_q0;
    end
  end

  assign Const_529 = (1'd0 ^ working_key[1053]);
  assign Const_530 = (1'd1 ^ working_key[1054]);
  assign Const_531 = (1'd0 ^ working_key[1055]);
  assign Const_532 = (1'd1 ^ working_key[1056]);
  assign Const_533 = (1'd1 ^ working_key[1057]);

  always @(*) begin
    if((((Const_529 == ap_CS_fsm_state49) | (Const_530 == ap_CS_fsm_state40) | (Const_531 == ap_CS_fsm_state46)) ^ working_key[1058]) == 1'b1) begin
      P_we0 = Const_532;
    end else begin
      P_we0 = Const_533;
    end
  end

  assign Const_534 = (1'd1 ^ working_key[1059]);
  assign Const_535 = (1'd1 ^ working_key[1060]);
  assign Const_536 = (1'd1 ^ working_key[1061]);
  assign Const_537 = (1'd1 ^ working_key[1062]);
  assign Const_538 = (1'd1 ^ working_key[1063]);

  always @(*) begin
    if((((Const_534 == ap_CS_fsm_state60) | (ap_start == Const_535) & (Const_536 == ap_CS_fsm_state1)) ^ working_key[1064]) == 1'b1) begin
      ap_done = Const_537;
    end else begin
      ap_done = Const_538;
    end
  end

  assign Const_539 = (1'd1 ^ working_key[1065]);
  assign Const_540 = (1'd1 ^ working_key[1066]);
  assign Const_541 = (1'd0 ^ working_key[1067]);
  assign Const_542 = (1'd0 ^ working_key[1068]);

  always @(*) begin
    if(((ap_start == Const_539) & (Const_540 == ap_CS_fsm_state1) ^ working_key[1069]) == 1'b1) begin
      ap_idle = Const_542;
    end else begin
      ap_idle = Const_541;
    end
  end

  assign Const_543 = (1'd0 ^ working_key[1070]);
  assign Const_544 = (1'd0 ^ working_key[1071]);
  assign Const_545 = (1'd0 ^ working_key[1072]);
  assign Const_546 = (1'd1 ^ working_key[1073]);
  assign Const_547 = (1'd1 ^ working_key[1074]);

  always @(*) begin
    if(((icmp_ln150_fu_2589_p2 == Const_543) & (icmp_ln147_reg_5407 == Const_544) & (icmp_ln204_reg_5387 == Const_545) & (icmp_ln178_reg_5248 == Const_546) & (Const_547 == ap_CS_fsm_state44) ^ working_key[1075]) == 1'b1) begin
      ap_phi_mux_p_0_i52_i_phi_fu_1041_p4 = p_0_i52_i_reg_1037;
    end else begin
      ap_phi_mux_p_0_i52_i_phi_fu_1041_p4 = div_0_i_i_reg_1015;
    end
  end

  assign Const_548 = (1'd0 ^ working_key[1076]);
  assign Const_549 = (1'd0 ^ working_key[1077]);
  assign Const_550 = (1'd0 ^ working_key[1078]);

  always @(*) begin
    if(((Const_548 == ap_CS_fsm_state60) ^ working_key[1079]) == 1'b1) begin
      ap_ready = Const_550;
    end else begin
      ap_ready = Const_549;
    end
  end

  assign Const_551 = (1'd1 ^ working_key[1080]);
  assign Const_552 = (1'd0 ^ working_key[1081]);

  always @(*) begin
    if(((Const_551 == ap_CS_fsm_state33) ^ working_key[1083]) == 1'b0) begin
      bitoff_address0 = zext_ln123_4_fu_2225_p1;
    end else if(((Const_552 == ap_CS_fsm_state2) ^ working_key[1082]) == 1'b1) begin
      bitoff_address0 = select_ln123_fu_1237_p3;
    end else begin
      bitoff_address0 = 'bx;
    end
  end

  assign Const_553 = (1'd1 ^ working_key[1084]);
  assign Const_554 = (1'd0 ^ working_key[1085]);

  always @(*) begin
    if(((Const_553 == ap_CS_fsm_state33) ^ working_key[1087]) == 1'b1) begin
      bitoff_address1 = zext_ln123_6_fu_2240_p1;
    end else if(((Const_554 == ap_CS_fsm_state2) ^ working_key[1086]) == 1'b1) begin
      bitoff_address1 = 'bx;
    end else begin
      bitoff_address1 = zext_ln123_1_fu_1256_p1;
    end
  end

  assign Const_555 = (1'd0 ^ working_key[1088]);
  assign Const_556 = (1'd1 ^ working_key[1089]);

  always @(*) begin
    if(((Const_555 == ap_CS_fsm_state33) ^ working_key[1091]) == 1'b1) begin
      bitoff_address2 = zext_ln123_8_fu_2255_p1;
    end else if(((Const_556 == ap_CS_fsm_state2) ^ working_key[1090]) == 1'b1) begin
      bitoff_address2 = 'bx;
    end else begin
      bitoff_address2 = zext_ln123_3_fu_1271_p1;
    end
  end

  assign Const_557 = (1'd1 ^ working_key[1092]);
  assign Const_558 = (1'd0 ^ working_key[1093]);
  assign Const_559 = (1'd1 ^ working_key[1094]);
  assign Const_560 = (1'd0 ^ working_key[1095]);

  always @(*) begin
    if((((Const_557 == ap_CS_fsm_state33) | (Const_558 == ap_CS_fsm_state2)) ^ working_key[1096]) == 1'b1) begin
      bitoff_ce0 = Const_560;
    end else begin
      bitoff_ce0 = Const_559;
    end
  end

  assign Const_561 = (1'd1 ^ working_key[1097]);
  assign Const_562 = (1'd0 ^ working_key[1098]);
  assign Const_563 = (1'd1 ^ working_key[1099]);
  assign Const_564 = (1'd1 ^ working_key[1100]);

  always @(*) begin
    if((((Const_561 == ap_CS_fsm_state33) | (Const_562 == ap_CS_fsm_state2)) ^ working_key[1101]) == 1'b1) begin
      bitoff_ce1 = Const_563;
    end else begin
      bitoff_ce1 = Const_564;
    end
  end

  assign Const_565 = (1'd0 ^ working_key[1102]);
  assign Const_566 = (1'd0 ^ working_key[1103]);
  assign Const_567 = (1'd1 ^ working_key[1104]);
  assign Const_568 = (1'd0 ^ working_key[1105]);

  always @(*) begin
    if((((Const_565 == ap_CS_fsm_state33) | (Const_566 == ap_CS_fsm_state2)) ^ working_key[1106]) == 1'b1) begin
      bitoff_ce2 = Const_568;
    end else begin
      bitoff_ce2 = Const_567;
    end
  end

  assign Const_569 = (1'd1 ^ working_key[1107]);
  assign Const_570 = (1'd0 ^ working_key[1108]);
  assign Const_571 = (1'd1 ^ working_key[1109]);

  always @(*) begin
    if(((Const_569 == ap_CS_fsm_state33) ^ working_key[1110]) == 1'b1) begin
      bitoff_ce3 = Const_571;
    end else begin
      bitoff_ce3 = Const_570;
    end
  end

  assign Const_572 = (1'd0 ^ working_key[1111]);
  assign Const_573 = (1'd0 ^ working_key[1112]);
  assign Const_574 = (1'd0 ^ working_key[1113]);

  always @(*) begin
    if(((Const_572 == ap_CS_fsm_state45) ^ working_key[1115]) == 1'b1) begin
      grp_fu_1093_p0 = temp_3_reg_5366;
    end else if((((Const_573 == ap_CS_fsm_state42) | (Const_574 == ap_CS_fsm_state48)) ^ working_key[1114]) == 1'b1) begin
      grp_fu_1093_p0 = 'bx;
    end else begin
      grp_fu_1093_p0 = P_q0;
    end
  end

  assign Const_575 = (1'd0 ^ working_key[1116]);
  assign Const_576 = (1'd1 ^ working_key[1117]);
  assign Const_577 = (1'd0 ^ working_key[1118]);
  assign Const_578 = (1'd1 ^ working_key[1119]);
  assign Const_579 = (1'd0 ^ working_key[1120]);
  assign Const_580 = (8'd83 ^ working_key[1128:1121]);
  assign Const_581 = (1'd0 ^ working_key[1129]);
  assign Const_582 = (8'd175 ^ working_key[1137:1130]);
  assign Const_583 = (1'd1 ^ working_key[1138]);
  assign Const_584 = (8'd7 ^ working_key[1146:1139]);
  assign Const_585 = (1'd0 ^ working_key[1147]);
  assign Const_586 = (8'd171 ^ working_key[1155:1148]);
  assign Const_587 = (1'd1 ^ working_key[1156]);
  assign Const_588 = (1'd0 ^ working_key[1157]);
  assign Const_589 = (1'd1 ^ working_key[1158]);
  assign Const_590 = (1'd1 ^ working_key[1159]);
  assign Const_591 = (8'd170 ^ working_key[1167:1160]);
  assign Const_592 = (1'd1 ^ working_key[1168]);
  assign Const_593 = (1'd0 ^ working_key[1169]);
  assign Const_594 = (1'd0 ^ working_key[1170]);
  assign Const_595 = (1'd0 ^ working_key[1171]);

  always @(*) begin
    if(((Const_575 == ap_CS_fsm_state24) ^ working_key[1183]) == 1'b0) begin
      s_address0 = sp_0_rec_i_cast_reg_5060;
    end else if(((Const_576 == ap_CS_fsm_state23) ^ working_key[1182]) == 1'b1) begin
      s_address0 = zext_ln146_fu_1959_p1;
    end else if(((Const_577 == ap_CS_fsm_state22) ^ working_key[1181]) == 1'b0) begin
      s_address0 = zext_ln144_fu_1911_p1;
    end else if(((Const_578 == ap_CS_fsm_state21) ^ working_key[1180]) == 1'b0) begin
      s_address0 = zext_ln142_fu_1877_p1;
    end else if(((Const_579 == ap_CS_fsm_state13) ^ working_key[1179]) == 1'b1) begin
      s_address0 = Const_580;
    end else if(((Const_581 == ap_CS_fsm_state12) ^ working_key[1178]) == 1'b0) begin
      s_address0 = Const_582;
    end else if(((Const_583 == ap_CS_fsm_state11) ^ working_key[1177]) == 1'b1) begin
      s_address0 = Const_584;
    end else if(((Const_585 == ap_CS_fsm_state10) ^ working_key[1176]) == 1'b0) begin
      s_address0 = Const_586;
    end else if(((Const_587 == ap_CS_fsm_state8) ^ working_key[1175]) == 1'b1) begin
      s_address0 = s_addr_2_reg_4709;
    end else if(((Const_588 == ap_CS_fsm_state6) & ((icmp_ln75_fu_1524_p2 == Const_589) | (Const_590 == and_ln72_reg_4687)) ^ working_key[1174]) == 1'b0) begin
      s_address0 = Const_591;
    end else if(((Const_592 == and_ln72_reg_4687) & (icmp_ln75_fu_1524_p2 == Const_593) & (Const_594 == ap_CS_fsm_state6) ^ working_key[1173]) == 1'b1) begin
      s_address0 = zext_ln76_1_fu_1536_p1;
    end else if(((Const_595 == ap_CS_fsm_state2) ^ working_key[1172]) == 1'b1) begin
      s_address0 = zext_ln60_fu_1138_p1;
    end else begin
      s_address0 = 'bx;
    end
  end

  assign Const_596 = (1'd1 ^ working_key[1184]);
  assign Const_597 = (1'd0 ^ working_key[1185]);
  assign Const_598 = (1'd1 ^ working_key[1186]);
  assign Const_599 = (1'd1 ^ working_key[1187]);
  assign Const_600 = (1'd0 ^ working_key[1188]);
  assign Const_601 = (1'd1 ^ working_key[1189]);
  assign Const_602 = (1'd1 ^ working_key[1190]);
  assign Const_603 = (1'd0 ^ working_key[1191]);
  assign Const_604 = (8'd108 ^ working_key[1199:1192]);
  assign Const_605 = (1'd1 ^ working_key[1200]);
  assign Const_606 = (8'd89 ^ working_key[1208:1201]);
  assign Const_607 = (1'd0 ^ working_key[1209]);
  assign Const_608 = (8'd89 ^ working_key[1217:1210]);

  always @(*) begin
    if(((Const_596 == ap_CS_fsm_state32) ^ working_key[1227]) == 1'b1) begin
      s_address1 = s_addr_19_reg_5235;
    end else if(((Const_597 == ap_CS_fsm_state31) ^ working_key[1226]) == 1'b0) begin
      s_address1 = p_0_rec_i_cast_fu_2078_p1;
    end else if(((Const_598 == ap_CS_fsm_state24) ^ working_key[1225]) == 1'b1) begin
      s_address1 = zext_ln138_fu_1964_p1;
    end else if(((Const_599 == ap_CS_fsm_state23) ^ working_key[1224]) == 1'b0) begin
      s_address1 = zext_ln145_fu_1948_p1;
    end else if(((Const_600 == ap_CS_fsm_state22) ^ working_key[1223]) == 1'b1) begin
      s_address1 = zext_ln143_fu_1900_p1;
    end else if(((Const_601 == ap_CS_fsm_state21) ^ working_key[1222]) == 1'b1) begin
      s_address1 = s_addr_10_reg_5065;
    end else if(((Const_602 == ap_CS_fsm_state20) ^ working_key[1221]) == 1'b0) begin
      s_address1 = zext_ln138_1_fu_1866_p1;
    end else if(((Const_603 == ap_CS_fsm_state13) ^ working_key[1220]) == 1'b1) begin
      s_address1 = Const_604;
    end else if(((Const_605 == ap_CS_fsm_state12) ^ working_key[1219]) == 1'b1) begin
      s_address1 = Const_606;
    end else if(((Const_607 == ap_CS_fsm_state11) ^ working_key[1218]) == 1'b1) begin
      s_address1 = 'bx;
    end else begin
      s_address1 = Const_608;
    end
  end

  assign Const_609 = (1'd0 ^ working_key[1228]);
  assign Const_610 = (1'd1 ^ working_key[1229]);
  assign Const_611 = (1'd0 ^ working_key[1230]);
  assign Const_612 = (1'd0 ^ working_key[1231]);
  assign Const_613 = (1'd1 ^ working_key[1232]);
  assign Const_614 = (1'd1 ^ working_key[1233]);
  assign Const_615 = (1'd0 ^ working_key[1234]);
  assign Const_616 = (1'd1 ^ working_key[1235]);
  assign Const_617 = (1'd0 ^ working_key[1236]);
  assign Const_618 = (1'd0 ^ working_key[1237]);
  assign Const_619 = (1'd0 ^ working_key[1238]);
  assign Const_620 = (1'd1 ^ working_key[1239]);
  assign Const_621 = (1'd0 ^ working_key[1240]);
  assign Const_622 = (1'd0 ^ working_key[1241]);
  assign Const_623 = (1'd0 ^ working_key[1242]);
  assign Const_624 = (1'd0 ^ working_key[1243]);
  assign Const_625 = (1'd0 ^ working_key[1244]);
  assign Const_626 = (1'd0 ^ working_key[1245]);

  always @(*) begin
    if((((Const_609 == ap_CS_fsm_state8) | (Const_610 == ap_CS_fsm_state12) | (Const_611 == ap_CS_fsm_state11) | (Const_612 == ap_CS_fsm_state10) | (Const_613 == ap_CS_fsm_state2) | (Const_614 == ap_CS_fsm_state24) | (Const_615 == ap_CS_fsm_state22) | (Const_616 == ap_CS_fsm_state23) | (Const_617 == ap_CS_fsm_state13) | (Const_618 == ap_CS_fsm_state21) | (Const_619 == and_ln72_reg_4687) & (icmp_ln75_fu_1524_p2 == Const_620) & (Const_621 == ap_CS_fsm_state6) | (Const_622 == ap_CS_fsm_state6) & ((icmp_ln75_fu_1524_p2 == Const_623) | (Const_624 == and_ln72_reg_4687))) ^ working_key[1246]) == 1'b1) begin
      s_ce0 = Const_626;
    end else begin
      s_ce0 = Const_625;
    end
  end

  assign Const_627 = (1'd1 ^ working_key[1247]);
  assign Const_628 = (1'd0 ^ working_key[1248]);
  assign Const_629 = (1'd1 ^ working_key[1249]);
  assign Const_630 = (1'd1 ^ working_key[1250]);
  assign Const_631 = (1'd0 ^ working_key[1251]);
  assign Const_632 = (1'd1 ^ working_key[1252]);
  assign Const_633 = (1'd0 ^ working_key[1253]);
  assign Const_634 = (1'd1 ^ working_key[1254]);
  assign Const_635 = (1'd0 ^ working_key[1255]);
  assign Const_636 = (1'd1 ^ working_key[1256]);
  assign Const_637 = (1'd0 ^ working_key[1257]);
  assign Const_638 = (1'd0 ^ working_key[1258]);

  always @(*) begin
    if((((Const_627 == ap_CS_fsm_state32) | (Const_628 == ap_CS_fsm_state31) | (Const_629 == ap_CS_fsm_state20) | (Const_630 == ap_CS_fsm_state12) | (Const_631 == ap_CS_fsm_state11) | (Const_632 == ap_CS_fsm_state24) | (Const_633 == ap_CS_fsm_state22) | (Const_634 == ap_CS_fsm_state23) | (Const_635 == ap_CS_fsm_state13) | (Const_636 == ap_CS_fsm_state21)) ^ working_key[1259]) == 1'b1) begin
      s_ce1 = Const_638;
    end else begin
      s_ce1 = Const_637;
    end
  end

  assign Const_639 = (1'd1 ^ working_key[1260]);
  assign Const_640 = (1'd0 ^ working_key[1261]);
  assign Const_641 = (1'd0 ^ working_key[1262]);

  always @(*) begin
    if(((Const_639 == ap_CS_fsm_state8) ^ working_key[1263]) == 1'b1) begin
      s_we0 = Const_641;
    end else begin
      s_we0 = Const_640;
    end
  end

  assign Const_642 = (1'd1 ^ working_key[1264]);
  assign Const_643 = (1'd0 ^ working_key[1265]);
  assign Const_644 = (1'd0 ^ working_key[1266]);

  always @(*) begin
    if(((Const_642 == ap_CS_fsm_state32) ^ working_key[1267]) == 1'b1) begin
      s_we1 = Const_644;
    end else begin
      s_we1 = Const_643;
    end
  end

  assign Const_645 = (1'd1 ^ working_key[1268]);
  assign Const_646 = (1'd0 ^ working_key[1269]);
  assign Const_647 = (1'd1 ^ working_key[1271]);
  assign Const_648 = (1'd1 ^ working_key[1272]);
  assign Const_649 = (1'd0 ^ working_key[1274]);
  assign Const_650 = (1'd0 ^ working_key[1275]);
  assign Const_651 = (1'd0 ^ working_key[1277]);
  assign Const_652 = (1'd1 ^ working_key[1278]);
  assign Const_653 = (1'd1 ^ working_key[1279]);
  assign Const_654 = (1'd1 ^ working_key[1281]);
  assign Const_655 = (1'd1 ^ working_key[1282]);
  assign Const_656 = (1'd1 ^ working_key[1284]);
  assign Const_657 = (1'd0 ^ working_key[1285]);
  assign Const_658 = (1'd0 ^ working_key[1287]);
  assign Const_659 = (1'd1 ^ working_key[1288]);
  assign Const_660 = (1'd1 ^ working_key[1290]);
  assign Const_661 = (1'd0 ^ working_key[1291]);
  assign Const_662 = (1'd0 ^ working_key[1292]);
  assign Const_663 = (1'd1 ^ working_key[1294]);
  assign Const_664 = (1'd0 ^ working_key[1295]);
  assign Const_665 = (1'd1 ^ working_key[1297]);
  assign Const_666 = (1'd0 ^ working_key[1298]);
  assign Const_667 = (1'd1 ^ working_key[1300]);
  assign Const_668 = (1'd0 ^ working_key[1301]);
  assign Const_669 = (1'd0 ^ working_key[1303]);
  assign Const_670 = (1'd0 ^ working_key[1304]);
  assign Const_671 = (1'd0 ^ working_key[1306]);
  assign Const_672 = (1'd1 ^ working_key[1307]);
  assign Const_673 = (1'd0 ^ working_key[1308]);
  assign Const_674 = (1'd0 ^ working_key[1309]);
  assign Const_675 = (1'd1 ^ working_key[1310]);
  assign Const_676 = (1'd0 ^ working_key[1311]);
  assign Const_677 = (1'd0 ^ working_key[1312]);
  assign Const_678 = (1'd0 ^ working_key[1313]);
  assign Const_679 = (1'd1 ^ working_key[1314]);
  assign Const_680 = (1'd0 ^ working_key[1315]);
  assign Const_681 = (1'd0 ^ working_key[1316]);
  assign Const_682 = (1'd1 ^ working_key[1317]);
  assign Const_683 = (1'd0 ^ working_key[1318]);
  assign Const_684 = (1'd1 ^ working_key[1319]);
  assign Const_685 = (1'd0 ^ working_key[1320]);
  assign Const_686 = (1'd0 ^ working_key[1321]);
  assign Const_687 = (1'd0 ^ working_key[1322]);
  assign Const_688 = (1'd1 ^ working_key[1323]);
  assign Const_689 = (1'd0 ^ working_key[1324]);
  assign Const_690 = (1'd1 ^ working_key[1327]);
  assign Const_691 = (1'd1 ^ working_key[1328]);
  assign Const_692 = (1'd1 ^ working_key[1330]);
  assign Const_693 = (1'd0 ^ working_key[1331]);
  assign Const_694 = (1'd0 ^ working_key[1333]);
  assign Const_695 = (1'd1 ^ working_key[1334]);

  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if(((ap_start == Const_645) & (Const_646 == ap_CS_fsm_state1) ^ working_key[1270]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if(((icmp_ln58_fu_1126_p2 == Const_647) & (Const_648 == ap_CS_fsm_state2) ^ working_key[1273]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end
      end
      ap_ST_fsm_state3: begin
        ap_NS_fsm = ap_ST_fsm_state2;
      end
      ap_ST_fsm_state4: begin
        if(((Const_649 == and_ln72_fu_1495_p2) & (Const_650 == ap_CS_fsm_state4) ^ working_key[1276]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end
      end
      ap_ST_fsm_state5: begin
        ap_NS_fsm = ap_ST_fsm_state6;
      end
      ap_ST_fsm_state6: begin
        if(((Const_651 == ap_CS_fsm_state6) & ((icmp_ln75_fu_1524_p2 == Const_652) | (Const_653 == and_ln72_reg_4687)) ^ working_key[1280]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state9;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end
      end
      ap_ST_fsm_state7: begin
        ap_NS_fsm = ap_ST_fsm_state8;
      end
      ap_ST_fsm_state8: begin
        ap_NS_fsm = ap_ST_fsm_state6;
      end
      ap_ST_fsm_state9: begin
        ap_NS_fsm = ap_ST_fsm_state10;
      end
      ap_ST_fsm_state10: begin
        if(((tmp_14_fu_1558_p3 == Const_654) & (Const_655 == ap_CS_fsm_state10) ^ working_key[1283]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state11;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state10;
        end
      end
      ap_ST_fsm_state11: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      ap_ST_fsm_state12: begin
        ap_NS_fsm = ap_ST_fsm_state13;
      end
      ap_ST_fsm_state13: begin
        ap_NS_fsm = ap_ST_fsm_state14;
      end
      ap_ST_fsm_state14: begin
        ap_NS_fsm = ap_ST_fsm_state15;
      end
      ap_ST_fsm_state15: begin
        ap_NS_fsm = ap_ST_fsm_state16;
      end
      ap_ST_fsm_state16: begin
        ap_NS_fsm = ap_ST_fsm_state17;
      end
      ap_ST_fsm_state17: begin
        ap_NS_fsm = ap_ST_fsm_state18;
      end
      ap_ST_fsm_state18: begin
        ap_NS_fsm = ap_ST_fsm_state19;
      end
      ap_ST_fsm_state19: begin
        ap_NS_fsm = ap_ST_fsm_state20;
      end
      ap_ST_fsm_state20: begin
        if(((icmp_ln135_fu_1848_p2 == Const_656) & (Const_657 == ap_CS_fsm_state20) ^ working_key[1286]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state29;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state21;
        end
      end
      ap_ST_fsm_state21: begin
        ap_NS_fsm = ap_ST_fsm_state22;
      end
      ap_ST_fsm_state22: begin
        ap_NS_fsm = ap_ST_fsm_state23;
      end
      ap_ST_fsm_state23: begin
        ap_NS_fsm = ap_ST_fsm_state24;
      end
      ap_ST_fsm_state24: begin
        ap_NS_fsm = ap_ST_fsm_state25;
      end
      ap_ST_fsm_state25: begin
        ap_NS_fsm = ap_ST_fsm_state26;
      end
      ap_ST_fsm_state26: begin
        ap_NS_fsm = ap_ST_fsm_state27;
      end
      ap_ST_fsm_state27: begin
        ap_NS_fsm = ap_ST_fsm_state28;
      end
      ap_ST_fsm_state28: begin
        ap_NS_fsm = ap_ST_fsm_state20;
      end
      ap_ST_fsm_state29: begin
        if(((tmp_15_fu_2052_p3 == Const_658) & (Const_659 == ap_CS_fsm_state29) ^ working_key[1289]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state30;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state31;
        end
      end
      ap_ST_fsm_state30: begin
        ap_NS_fsm = ap_ST_fsm_state29;
      end
      ap_ST_fsm_state31: begin
        if(((Const_660 == ap_CS_fsm_state31) & ((icmp_ln158_fu_2083_p2 == Const_661) | (icmp_ln72_reg_4683 == Const_662)) ^ working_key[1293]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state32;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state33;
        end
      end
      ap_ST_fsm_state32: begin
        ap_NS_fsm = ap_ST_fsm_state31;
      end
      ap_ST_fsm_state33: begin
        if(((icmp_ln178_fu_2101_p2 == Const_663) & (Const_664 == ap_CS_fsm_state33) ^ working_key[1296]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state50;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state34;
        end
      end
      ap_ST_fsm_state34: begin
        ap_NS_fsm = ap_ST_fsm_state35;
      end
      ap_ST_fsm_state35: begin
        if(((icmp_ln186_fu_2443_p2 == Const_665) & (Const_666 == ap_CS_fsm_state35) ^ working_key[1299]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state36;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state37;
        end
      end
      ap_ST_fsm_state36: begin
        ap_NS_fsm = ap_ST_fsm_state35;
      end
      ap_ST_fsm_state37: begin
        if(((icmp_ln192_fu_2480_p2 == Const_667) & (Const_668 == ap_CS_fsm_state37) ^ working_key[1302]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state38;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state39;
        end
      end
      ap_ST_fsm_state38: begin
        ap_NS_fsm = ap_ST_fsm_state37;
      end
      ap_ST_fsm_state39: begin
        if(((icmp_ln194_fu_2497_p2 == Const_669) & (Const_670 == ap_CS_fsm_state39) ^ working_key[1305]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state41;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state40;
        end
      end
      ap_ST_fsm_state40: begin
        ap_NS_fsm = ap_ST_fsm_state39;
      end
      ap_ST_fsm_state41: begin
        ap_NS_fsm = ap_ST_fsm_state42;
      end
      ap_ST_fsm_state42: begin
        ap_NS_fsm = ap_ST_fsm_state43;
      end
      ap_ST_fsm_state43: begin
        ap_NS_fsm = ap_ST_fsm_state44;
      end
      ap_ST_fsm_state44: begin
        if(((Const_671 == ap_CS_fsm_state44) & ((icmp_ln178_reg_5248 == Const_672) | ((icmp_ln206_fu_2677_p2 == Const_673) & (icmp_ln204_reg_5387 == Const_674) | (icmp_ln215_fu_2657_p2 == Const_675) & (icmp_ln150_fu_2589_p2 == Const_676) & (icmp_ln204_reg_5387 == Const_677) | (icmp_ln215_fu_2657_p2 == Const_678) & (icmp_ln147_reg_5407 == Const_679) & (icmp_ln204_reg_5387 == Const_680))) ^ working_key[1326]) == 1'b0) begin
          ap_NS_fsm = ap_ST_fsm_state51;
        end else if(((Const_681 == ap_CS_fsm_state44) & ((icmp_ln147_reg_5407 == Const_682) & (icmp_ln215_fu_2657_p2 == Const_683) & (icmp_ln204_reg_5387 == Const_684) & (icmp_ln178_reg_5248 == Const_685) | (icmp_ln150_fu_2589_p2 == Const_686) & (icmp_ln215_fu_2657_p2 == Const_687) & (icmp_ln204_reg_5387 == Const_688) & (icmp_ln178_reg_5248 == Const_689)) ^ working_key[1325]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state44;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state45;
        end
      end
      ap_ST_fsm_state45: begin
        ap_NS_fsm = ap_ST_fsm_state46;
      end
      ap_ST_fsm_state46: begin
        ap_NS_fsm = ap_ST_fsm_state47;
      end
      ap_ST_fsm_state47: begin
        if(((icmp_ln223_fu_2788_p2 == Const_690) & (Const_691 == ap_CS_fsm_state47) ^ working_key[1329]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state48;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state41;
        end
      end
      ap_ST_fsm_state48: begin
        ap_NS_fsm = ap_ST_fsm_state49;
      end
      ap_ST_fsm_state49: begin
        ap_NS_fsm = ap_ST_fsm_state47;
      end
      ap_ST_fsm_state50: begin
        if(((icmp_ln180_fu_3008_p2 == Const_692) & (Const_693 == ap_CS_fsm_state50) ^ working_key[1332]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state50;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state44;
        end
      end
      ap_ST_fsm_state51: begin
        if(((icmp_ln253_fu_3025_p2 == Const_694) & (Const_695 == ap_CS_fsm_state51) ^ working_key[1335]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state52;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state54;
        end
      end
      ap_ST_fsm_state52: begin
        ap_NS_fsm = ap_ST_fsm_state53;
      end
      ap_ST_fsm_state53: begin
        ap_NS_fsm = ap_ST_fsm_state51;
      end
      ap_ST_fsm_state54: begin
        ap_NS_fsm = ap_ST_fsm_state55;
      end
      ap_ST_fsm_state55: begin
        ap_NS_fsm = ap_ST_fsm_state56;
      end
      ap_ST_fsm_state56: begin
        ap_NS_fsm = ap_ST_fsm_state57;
      end
      ap_ST_fsm_state57: begin
        ap_NS_fsm = ap_ST_fsm_state58;
      end
      ap_ST_fsm_state58: begin
        ap_NS_fsm = ap_ST_fsm_state59;
      end
      ap_ST_fsm_state59: begin
        ap_NS_fsm = ap_ST_fsm_state60;
      end
      ap_ST_fsm_state60: begin
        ap_NS_fsm = ap_ST_fsm_state1;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign ACF_d0 = { { shl_ln187_fu_2464_p2[31:16] } };
  assign Const_696 = (3'd4 ^ working_key[1338:1336]);
  assign LARc_addr_10_reg_5633 = Const_696;
  assign Const_697 = (3'd2 ^ working_key[1341:1339]);
  assign LARc_addr_11_reg_5638 = Const_697;
  assign Const_698 = (3'd7 ^ working_key[1344:1342]);
  assign LARc_addr_6_reg_5577 = Const_698;
  assign Const_699 = (3'd1 ^ working_key[1347:1345]);
  assign LARc_addr_7_reg_5582 = Const_699;
  assign Const_700 = (3'd6 ^ working_key[1350:1348]);
  assign LARc_addr_8_reg_5607 = Const_700;
  assign Const_701 = (3'd7 ^ working_key[1353:1351]);
  assign LARc_addr_9_reg_5612 = Const_701;
  assign Const_702 = (4'd4 ^ working_key[1357:1354]);
  assign L_ACF_addr_1_reg_4748 = Const_702;
  assign Const_703 = (4'd1 ^ working_key[1361:1358]);
  assign L_ACF_addr_2_reg_4776 = Const_703;
  assign Const_704 = (4'd14 ^ working_key[1365:1362]);
  assign L_ACF_addr_3_reg_4782 = Const_704;
  assign Const_705 = (4'd11 ^ working_key[1369:1366]);
  assign L_ACF_addr_4_reg_4885 = Const_705;
  assign Const_706 = (4'd0 ^ working_key[1373:1370]);
  assign L_ACF_addr_5_reg_4911 = Const_706;
  assign Const_707 = (4'd3 ^ working_key[1377:1374]);
  assign L_ACF_addr_6_reg_4967 = Const_707;
  assign Const_708 = (4'd13 ^ working_key[1381:1378]);
  assign L_ACF_addr_7_reg_5023 = Const_708;
  assign Const_709 = (64'd5392271837434522283 ^ working_key[1445:1382]);
  assign L_num_1_fu_2595_p2 = (working_key[1446] == 1'b1)? L_num_0_i_i_reg_1006 >> Const_709 : L_num_0_i_i_reg_1006 << Const_709;
  assign L_num_2_fu_2606_p2 = (working_key[1447] == 1'b1)? L_num_1_fu_2595_p2 - sext_ln139_reg_5396 : L_num_1_fu_2595_p2 * sext_ln139_reg_5396;
  assign Const_710 = (1'd1 ^ working_key[1448]);
  assign L_num_3_fu_2611_p3 = ((((working_key[1449] == 1'b1)? icmp_ln155_fu_2601_p2[0:0] === Const_710 : icmp_ln155_fu_2601_p2[0:0] == Const_710) ^ working_key[1450]) == 1'b1)? L_num_1_fu_2595_p2 : L_num_2_fu_2606_p2;
  assign a_assign_1_fu_1143_p3 = { { smax_0_i_reg_839 }, { 16'd0 } };
  assign Const_711 = (4'd2 ^ working_key[1454:1451]);
  assign add_ln123_1_fu_1362_p2 = (working_key[1455] == 1'b1)? Const_711 - bitoff_q2 : Const_711 + bitoff_q2;
  assign Const_712 = (5'd13 ^ working_key[1460:1456]);
  assign add_ln123_2_fu_2371_p2 = (working_key[1461] == 1'b1)? Const_712 + zext_ln123_5_fu_2367_p1 : Const_712 << zext_ln123_5_fu_2367_p1;
  assign Const_713 = (5'd5 ^ working_key[1466:1462]);
  assign add_ln123_3_fu_2381_p2 = (working_key[1467] == 1'b1)? Const_713 + zext_ln123_7_fu_2377_p1 : Const_713 << zext_ln123_7_fu_2377_p1;
  assign Const_714 = (4'd1 ^ working_key[1471:1468]);
  assign add_ln123_4_fu_2387_p2 = (working_key[1472] == 1'b1)? Const_714 + bitoff_q2 : Const_714 * bitoff_q2;
  assign Const_715 = (4'd13 ^ working_key[1476:1473]);
  assign add_ln123_5_fu_2397_p2 = (working_key[1477] == 1'b1)? Const_715 + bitoff_q3 : Const_715 >> bitoff_q3;
  assign Const_716 = (4'd3 ^ working_key[1481:1478]);
  assign add_ln123_fu_1352_p2 = (working_key[1482] == 1'b1)? Const_716 + bitoff_q1 : Const_716 - bitoff_q1;
  assign add_ln126_1_fu_1757_p2 = (working_key[1483] == 1'b1)? reg_1104 - sext_ln111_2_fu_1754_p1 : reg_1104 + sext_ln111_2_fu_1754_p1;
  assign add_ln126_3_fu_1766_p2 = (working_key[1484] == 1'b1)? sext_ln126_3_fu_1763_p1 + add_ln126_1_fu_1757_p2 : sext_ln126_3_fu_1763_p1 >> add_ln126_1_fu_1757_p2;
  assign add_ln126_7_fu_1672_p2 = (working_key[1485] == 1'b1)? sext_ln126_5_fu_1669_p1 >> sext_ln126_4_fu_1666_p1 : sext_ln126_5_fu_1669_p1 + sext_ln126_4_fu_1666_p1;
  assign add_ln126_fu_1775_p2 = (working_key[1486] == 1'b1)? sext_ln126_6_fu_1772_p1 + add_ln126_3_fu_1766_p2 : sext_ln126_6_fu_1772_p1 << add_ln126_3_fu_1766_p2;
  assign add_ln127_1_fu_1678_p2 = (working_key[1487] == 1'b1)? reg_1109 + sext_ln94_fu_1623_p1 : reg_1109 >> sext_ln94_fu_1623_p1;
  assign add_ln127_3_fu_1687_p2 = (working_key[1488] == 1'b1)? sext_ln127_1_fu_1684_p1 - add_ln127_1_fu_1678_p2 : sext_ln127_1_fu_1684_p1 + add_ln127_1_fu_1678_p2;
  assign add_ln127_fu_1699_p2 = (working_key[1489] == 1'b1)? sext_ln127_6_fu_1696_p1 - add_ln127_3_fu_1687_p2 : sext_ln127_6_fu_1696_p1 + add_ln127_3_fu_1687_p2;
  assign add_ln128_2_fu_1708_p2 = (working_key[1490] == 1'b1)? sext_ln128_1_fu_1705_p1 + reg_1114 : sext_ln128_1_fu_1705_p1 - reg_1114;
  assign add_ln128_5_fu_1720_p2 = (working_key[1491] == 1'b1)? sext_ln128_3_fu_1717_p1 << sext_ln128_2_fu_1714_p1 : sext_ln128_3_fu_1717_p1 + sext_ln128_2_fu_1714_p1;
  assign add_ln128_fu_1730_p2 = (working_key[1492] == 1'b1)? sext_ln128_4_fu_1726_p1 + add_ln128_2_fu_1708_p2 : sext_ln128_4_fu_1726_p1 - add_ln128_2_fu_1708_p2;
  assign add_ln129_2_fu_1785_p2 = (working_key[1493] == 1'b1)? sext_ln129_1_fu_1782_p1 + reg_1118 : sext_ln129_1_fu_1782_p1 << reg_1118;
  assign add_ln129_fu_1794_p2 = (working_key[1494] == 1'b1)? sext_ln129_2_fu_1791_p1 + add_ln129_2_fu_1785_p2 : sext_ln129_2_fu_1791_p1 >> add_ln129_2_fu_1785_p2;
  assign add_ln130_1_fu_1800_p2 = (working_key[1495] == 1'b1)? reg_1109 + sext_ln109_fu_1751_p1 : reg_1109 - sext_ln109_fu_1751_p1;
  assign add_ln130_fu_1809_p2 = (working_key[1496] == 1'b1)? sext_ln130_1_fu_1806_p1 + add_ln130_1_fu_1800_p2 : sext_ln130_1_fu_1806_p1 - add_ln130_1_fu_1800_p2;
  assign add_ln131_1_fu_1736_p2 = (working_key[1497] == 1'b1)? L_ACF_q0 + sext_ln116_fu_1641_p1 : L_ACF_q0 >> sext_ln116_fu_1641_p1;
  assign add_ln131_fu_1745_p2 = (working_key[1498] == 1'b1)? sext_ln131_1_fu_1742_p1 + add_ln131_1_fu_1736_p2 : sext_ln131_1_fu_1742_p1 * add_ln131_1_fu_1736_p2;
  assign add_ln132_fu_1818_p2 = (working_key[1499] == 1'b1)? sext_ln132_1_fu_1815_p1 >> L_ACF_q1 : sext_ln132_1_fu_1815_p1 + L_ACF_q1;
  assign add_ln133_fu_1827_p2 = (working_key[1500] == 1'b1)? L_ACF_q0 + sext_ln133_fu_1824_p1 : L_ACF_q0 - sext_ln133_fu_1824_p1;
  assign Const_717 = (8'd66 ^ working_key[1508:1501]);
  assign add_ln138_1_fu_1860_p2 = (working_key[1509] == 1'b1)? sp_0_rec_i_reg_894 + Const_717 : sp_0_rec_i_reg_894 >> Const_717;
  assign Const_718 = (8'd171 ^ working_key[1517:1510]);
  assign add_ln138_fu_1854_p2 = (working_key[1518] == 1'b1)? sp_0_rec_i_reg_894 - Const_718 : sp_0_rec_i_reg_894 + Const_718;
  assign add_ln140_fu_1971_p2 = (working_key[1519] == 1'b1)? sext_ln140_1_fu_1968_p1 + empty_57_reg_884 : sext_ln140_1_fu_1968_p1 - empty_57_reg_884;
  assign add_ln141_fu_1919_p2 = (working_key[1520] == 1'b1)? reg_1104 << sext_ln141_1_fu_1916_p1 : reg_1104 + sext_ln141_1_fu_1916_p1;
  assign add_ln142_1_fu_1928_p2 = (working_key[1521] == 1'b1)? reg_1109 + sext_ln142_1_fu_1925_p1 : reg_1109 - sext_ln142_1_fu_1925_p1;
  assign Const_719 = (8'd12 ^ working_key[1529:1522]);
  assign add_ln142_fu_1871_p2 = (working_key[1530] == 1'b1)? sp_0_rec_i_reg_894 >> Const_719 : sp_0_rec_i_reg_894 + Const_719;
  assign add_ln143_1_fu_1981_p2 = (working_key[1531] == 1'b1)? reg_1114 + sext_ln143_1_fu_1978_p1 : reg_1114 >> sext_ln143_1_fu_1978_p1;
  assign Const_720 = (8'd175 ^ working_key[1539:1532]);
  assign add_ln143_fu_1894_p2 = (working_key[1540] == 1'b1)? sp_0_rec_i_reg_894 - Const_720 : sp_0_rec_i_reg_894 + Const_720;
  assign add_ln144_1_fu_1990_p2 = (working_key[1541] == 1'b1)? reg_1118 + sext_ln144_1_fu_1987_p1 : reg_1118 << sext_ln144_1_fu_1987_p1;
  assign Const_721 = (8'd174 ^ working_key[1549:1542]);
  assign add_ln144_fu_1905_p2 = (working_key[1550] == 1'b1)? sp_0_rec_i_reg_894 * Const_721 : sp_0_rec_i_reg_894 + Const_721;
  assign add_ln145_1_fu_2007_p2 = (working_key[1551] == 1'b1)? reg_1104 + sext_ln145_1_fu_2004_p1 : reg_1104 * sext_ln145_1_fu_2004_p1;
  assign Const_722 = (8'd239 ^ working_key[1559:1552]);
  assign add_ln145_fu_1942_p2 = (working_key[1560] == 1'b1)? sp_0_rec_i_reg_894 + Const_722 : sp_0_rec_i_reg_894 << Const_722;
  assign add_ln146_1_fu_2016_p2 = (working_key[1561] == 1'b1)? reg_1109 >> sext_ln146_1_fu_2013_p1 : reg_1109 + sext_ln146_1_fu_2013_p1;
  assign Const_723 = (8'd175 ^ working_key[1569:1562]);
  assign add_ln146_fu_1953_p2 = (working_key[1570] == 1'b1)? sp_0_rec_i_reg_894 << Const_723 : sp_0_rec_i_reg_894 + Const_723;
  assign add_ln147_fu_2033_p2 = (working_key[1571] == 1'b1)? reg_1114 * sext_ln147_1_fu_2030_p1 : reg_1114 + sext_ln147_1_fu_2030_p1;
  assign add_ln148_fu_2042_p2 = (working_key[1572] == 1'b1)? reg_1118 + sext_ln148_1_fu_2039_p1 : reg_1118 << sext_ln148_1_fu_2039_p1;
  assign Const_724 = (4'd11 ^ working_key[1576:1573]);
  assign add_ln150_fu_2583_p2 = (working_key[1577] == 1'b1)? k_0_i_i_reg_1026 + Const_724 : k_0_i_i_reg_1026 * Const_724;
  assign Const_725 = (8'd155 ^ working_key[1585:1578]);
  assign add_ln159_fu_2089_p2 = (working_key[1586] == 1'b1)? p_0_rec_i_reg_917 * Const_725 : p_0_rec_i_reg_917 + Const_725;
  assign Const_726 = (4'd6 ^ working_key[1590:1587]);
  assign add_ln181_fu_3014_p2 = (working_key[1591] == 1'b1)? p_0_rec_i1_reg_1071 + Const_726 : p_0_rec_i1_reg_1071 << Const_726;
  assign Const_727 = (32'd187357845 ^ working_key[1623:1592]);
  assign add_ln199_2_fu_2815_p2 = (working_key[1624] == 1'b1)? indvars_iv142_reg_961 + Const_727 : indvars_iv142_reg_961 >> Const_727;
  assign Const_728 = (4'd10 ^ working_key[1628:1625]);
  assign add_ln199_fu_2527_p2 = (working_key[1629] == 1'b1)? p_1_rec_i_reg_985 * Const_728 : p_1_rec_i_reg_985 + Const_728;
  assign Const_729 = (32'd2695539364 ^ working_key[1661:1630]);
  assign add_ln207_fu_2683_p2 = (working_key[1662] == 1'b1)? Const_729 * p_2_rec_i_reg_1049 : Const_729 + p_2_rec_i_reg_1049;
  assign Const_730 = (4'd4 ^ working_key[1666:1663]);
  assign add_ln253_fu_3031_p2 = (working_key[1667] == 1'b1)? p_0_rec_i16_reg_1082 + Const_730 : p_0_rec_i16_reg_1082 * Const_730;
  assign Const_731 = (8'd138 ^ working_key[1675:1668]);
  assign add_ln304_fu_3634_p2 = (working_key[1676] == 1'b1)? sext_ln304_fu_3608_p1 >> Const_731 : sext_ln304_fu_3608_p1 + Const_731;
  assign Const_732 = (8'd69 ^ working_key[1684:1677]);
  assign add_ln305_fu_3699_p2 = (working_key[1685] == 1'b1)? sext_ln305_fu_3673_p1 * Const_732 : sext_ln305_fu_3673_p1 + Const_732;
  assign Const_733 = (8'd197 ^ working_key[1693:1686]);
  assign add_ln306_fu_3870_p2 = (working_key[1694] == 1'b1)? sext_ln306_fu_3844_p1 << Const_733 : sext_ln306_fu_3844_p1 + Const_733;
  assign Const_734 = (8'd53 ^ working_key[1702:1695]);
  assign add_ln307_fu_3935_p2 = (working_key[1703] == 1'b1)? sext_ln307_fu_3909_p1 + Const_734 : sext_ln307_fu_3909_p1 << Const_734;
  assign Const_735 = (8'd98 ^ working_key[1711:1704]);
  assign add_ln309_fu_4060_p2 = (working_key[1712] == 1'b1)? sext_ln309_fu_4034_p1 << Const_735 : sext_ln309_fu_4034_p1 + Const_735;
  assign Const_736 = (8'd85 ^ working_key[1720:1713]);
  assign add_ln310_fu_4125_p2 = (working_key[1721] == 1'b1)? sext_ln310_fu_4099_p1 + Const_736 : sext_ln310_fu_4099_p1 >> Const_736;
  assign Const_737 = (8'd94 ^ working_key[1729:1722]);
  assign add_ln311_fu_4190_p2 = (working_key[1730] == 1'b1)? sext_ln311_fu_4164_p1 + Const_737 : sext_ln311_fu_4164_p1 >> Const_737;
  assign Const_738 = (8'd160 ^ working_key[1738:1731]);
  assign add_ln312_fu_4255_p2 = (working_key[1739] == 1'b1)? sext_ln312_fu_4229_p1 - Const_738 : sext_ln312_fu_4229_p1 + Const_738;
  assign add_ln40_10_fu_2976_p2 = (working_key[1740] == 1'b1)? temp_7_reg_5518 + K_load_reg_5506 : temp_7_reg_5518 >> K_load_reg_5506;
  assign Const_739 = (16'd16397 ^ working_key[1756:1741]);
  assign add_ln40_11_fu_3983_p2 = (working_key[1757] == 1'b1)? temp_16_reg_5653 << Const_739 : temp_16_reg_5653 + Const_739;
  assign Const_740 = (16'd22061 ^ working_key[1773:1758]);
  assign add_ln40_12_fu_4013_p2 = (working_key[1774] == 1'b1)? temp_17_reg_5659 >> Const_740 : temp_17_reg_5659 + Const_740;
  assign add_ln40_1_fu_2754_p2 = (working_key[1775] == 1'b1)? temp_5_fu_2715_p3 + reg_1122 : temp_5_fu_2715_p3 >> reg_1122;
  assign Const_741 = (16'd43306 ^ working_key[1791:1776]);
  assign add_ln40_2_fu_3307_p2 = (working_key[1792] == 1'b1)? temp_9_fu_3271_p4 - Const_741 : temp_9_fu_3271_p4 + Const_741;
  assign Const_742 = (16'd23893 ^ working_key[1808:1793]);
  assign add_ln40_3_fu_3389_p2 = (working_key[1809] == 1'b1)? temp_10_fu_3353_p4 * Const_742 : temp_10_fu_3353_p4 + Const_742;
  assign Const_743 = (16'd44155 ^ working_key[1825:1810]);
  assign add_ln40_4_fu_3429_p2 = (working_key[1826] == 1'b1)? temp_11_fu_3395_p3 * Const_743 : temp_11_fu_3395_p3 + Const_743;
  assign Const_744 = (16'd47698 ^ working_key[1842:1827]);
  assign add_ln40_5_fu_3501_p2 = (working_key[1843] == 1'b1)? temp_12_fu_3475_p4 + Const_744 : temp_12_fu_3475_p4 * Const_744;
  assign add_ln40_6_fu_2917_p2 = (working_key[1844] == 1'b1)? temp_6_reg_5512 + reg_1122 : temp_6_reg_5512 * reg_1122;
  assign Const_745 = (16'd11019 ^ working_key[1860:1845]);
  assign add_ln40_7_fu_3757_p2 = (working_key[1861] == 1'b1)? temp_13_reg_5617 + Const_745 : temp_13_reg_5617 - Const_745;
  assign Const_746 = (16'd53844 ^ working_key[1877:1862]);
  assign add_ln40_8_fu_3796_p2 = (working_key[1878] == 1'b1)? temp_14_fu_3762_p3 + Const_746 : temp_14_fu_3762_p3 - Const_746;
  assign Const_747 = (16'd43183 ^ working_key[1894:1879]);
  assign add_ln40_9_fu_3586_p2 = (working_key[1895] == 1'b1)? temp_15_fu_3560_p4 + Const_747 : temp_15_fu_3560_p4 * Const_747;
  assign Const_748 = (16'd11178 ^ working_key[1911:1896]);
  assign add_ln40_fu_3225_p2 = (working_key[1912] == 1'b1)? temp_8_fu_3189_p4 << Const_748 : temp_8_fu_3189_p4 + Const_748;
  assign add_ln50_1_fu_3265_p2 = (working_key[1913] == 1'b1)? sext_ln50_3_fu_3261_p1 << sext_ln50_2_fu_3249_p1 : sext_ln50_3_fu_3261_p1 + sext_ln50_2_fu_3249_p1;
  assign add_ln50_2_fu_3347_p2 = (working_key[1914] == 1'b1)? sext_ln50_5_fu_3343_p1 - sext_ln50_4_fu_3331_p1 : sext_ln50_5_fu_3343_p1 + sext_ln50_4_fu_3331_p1;
  assign add_ln50_3_fu_3469_p2 = (working_key[1915] == 1'b1)? sext_ln50_7_fu_3465_p1 + sext_ln50_6_fu_3453_p1 : sext_ln50_7_fu_3465_p1 - sext_ln50_6_fu_3453_p1;
  assign add_ln50_fu_3183_p2 = (working_key[1916] == 1'b1)? sext_ln50_1_fu_3179_p1 - sext_ln50_fu_3167_p1 : sext_ln50_1_fu_3179_p1 + sext_ln50_fu_3167_p1;
  assign Const_749 = (3'd2 ^ working_key[1919:1917]);
  assign add_ln76_fu_1505_p2 = (working_key[1920] == 1'b1)? Const_749 << trunc_ln76_reg_4691 : Const_749 + trunc_ln76_reg_4691;
  assign and_ln263_fu_3131_p2 = (working_key[1921] == 1'b1)? xor_ln259_fu_3125_p2 & icmp_ln263_fu_3093_p2 : xor_ln259_fu_3125_p2 | icmp_ln263_fu_3093_p2;
  assign and_ln58_1_fu_2827_p2 = (working_key[1922] == 1'b1)? icmp_ln58_3_fu_2821_p2 | icmp_ln58_1_reg_5451 : icmp_ln58_3_fu_2821_p2 & icmp_ln58_1_reg_5451;
  assign and_ln58_2_fu_2857_p2 = (working_key[1923] == 1'b1)? icmp_ln58_1_reg_5451 & grp_fu_1093_p2 : icmp_ln58_1_reg_5451 << grp_fu_1093_p2;
  assign and_ln58_fu_2694_p2 = (working_key[1924] == 1'b1)? icmp_ln58_1_fu_2689_p2 << grp_fu_1093_p2 : icmp_ln58_1_fu_2689_p2 & grp_fu_1093_p2;
  assign and_ln72_fu_1495_p2 = (working_key[1925] == 1'b1)? icmp_ln72_fu_1483_p2 & icmp_ln72_2_fu_1489_p2 : icmp_ln72_fu_1483_p2 << icmp_ln72_2_fu_1489_p2;
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];
  assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];
  assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];
  assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];
  assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];
  assign ap_CS_fsm_state21 = ap_CS_fsm[32'd20];
  assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];
  assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];
  assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];
  assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];
  assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];
  assign ap_CS_fsm_state27 = ap_CS_fsm[32'd26];
  assign ap_CS_fsm_state28 = ap_CS_fsm[32'd27];
  assign ap_CS_fsm_state29 = ap_CS_fsm[32'd28];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state30 = ap_CS_fsm[32'd29];
  assign ap_CS_fsm_state31 = ap_CS_fsm[32'd30];
  assign ap_CS_fsm_state32 = ap_CS_fsm[32'd31];
  assign ap_CS_fsm_state33 = ap_CS_fsm[32'd32];
  assign ap_CS_fsm_state34 = ap_CS_fsm[32'd33];
  assign ap_CS_fsm_state35 = ap_CS_fsm[32'd34];
  assign ap_CS_fsm_state36 = ap_CS_fsm[32'd35];
  assign ap_CS_fsm_state37 = ap_CS_fsm[32'd36];
  assign ap_CS_fsm_state38 = ap_CS_fsm[32'd37];
  assign ap_CS_fsm_state39 = ap_CS_fsm[32'd38];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state40 = ap_CS_fsm[32'd39];
  assign ap_CS_fsm_state41 = ap_CS_fsm[32'd40];
  assign ap_CS_fsm_state42 = ap_CS_fsm[32'd41];
  assign ap_CS_fsm_state43 = ap_CS_fsm[32'd42];
  assign ap_CS_fsm_state44 = ap_CS_fsm[32'd43];
  assign ap_CS_fsm_state45 = ap_CS_fsm[32'd44];
  assign ap_CS_fsm_state46 = ap_CS_fsm[32'd45];
  assign ap_CS_fsm_state47 = ap_CS_fsm[32'd46];
  assign ap_CS_fsm_state48 = ap_CS_fsm[32'd47];
  assign ap_CS_fsm_state49 = ap_CS_fsm[32'd48];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state50 = ap_CS_fsm[32'd49];
  assign ap_CS_fsm_state51 = ap_CS_fsm[32'd50];
  assign ap_CS_fsm_state52 = ap_CS_fsm[32'd51];
  assign ap_CS_fsm_state53 = ap_CS_fsm[32'd52];
  assign ap_CS_fsm_state54 = ap_CS_fsm[32'd53];
  assign ap_CS_fsm_state55 = ap_CS_fsm[32'd54];
  assign ap_CS_fsm_state56 = ap_CS_fsm[32'd55];
  assign ap_CS_fsm_state57 = ap_CS_fsm[32'd56];
  assign ap_CS_fsm_state58 = ap_CS_fsm[32'd57];
  assign ap_CS_fsm_state59 = ap_CS_fsm[32'd58];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state60 = ap_CS_fsm[32'd59];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign bitoff_address3 = zext_ln123_10_fu_2270_p1;
  assign div_fu_2629_p3 = { { trunc_ln155_fu_2625_p1 }, { xor_ln155_fu_2619_p2 } };
  assign empty_65_fu_2663_p1 = p_2_rec_i_reg_1049[4:0];
  assign Const_750 = (16'd45738 ^ working_key[1941:1926]);
  assign Const_751 = (1'd1 ^ working_key[1943]);
  assign Const_752 = (1'd1 ^ working_key[1944]);
  assign grp_fu_1093_p2 = ((((working_key[1942] == 1'b1)? grp_fu_1093_p0 == Const_750 : grp_fu_1093_p0 === Const_750) ^ working_key[1945]) == 1'b1)? Const_751 : Const_752;
  assign grp_fu_4288_p0 = zext_ln75_reg_4696;
  assign Const_753 = (16'd58541 ^ working_key[1961:1946]);
  assign grp_fu_4288_p2 = Const_753;
  assign grp_fu_4390_p0 = sext_ln91_reg_4810;
  assign grp_fu_4390_p1 = sext_ln91_reg_4810;
  assign grp_fu_4397_p0 = sext_ln96_1_reg_4836;
  assign grp_fu_4397_p1 = sext_ln96_1_reg_4836;
  assign grp_fu_4403_p0 = sext_ln100_1_reg_4854;
  assign grp_fu_4403_p1 = sext_ln93_1_reg_4818;
  assign grp_fu_4410_p0 = sext_ln105_1_reg_4871;
  assign grp_fu_4410_p1 = sext_ln105_1_reg_4871;
  assign grp_fu_4416_p0 = sext_ln105_1_reg_4871;
  assign grp_fu_4416_p1 = sext_ln93_1_reg_4818;
  assign grp_fu_4430_p0 = sext_ln111_1_reg_4896;
  assign grp_fu_4430_p1 = sext_ln100_1_reg_4854;
  assign grp_fu_4437_p0 = sext_ln111_1_reg_4896;
  assign grp_fu_4437_p1 = sext_ln96_1_reg_4836;
  assign grp_fu_4442_p0 = sext_ln111_1_reg_4896;
  assign grp_fu_4442_p1 = sext_ln93_1_reg_4818;
  assign grp_fu_4447_p0 = sext_ln126_1_fu_1662_p1;
  assign grp_fu_4447_p1 = sext_ln126_1_fu_1662_p1;
  assign grp_fu_4456_p0 = sext_ln100_reg_4849;
  assign grp_fu_4456_p1 = sext_ln111_reg_4891;
  assign grp_fu_4465_p0 = sext_ln126_1_fu_1662_p1;
  assign grp_fu_4465_p1 = sext_ln111_1_reg_4896;
  assign grp_fu_4473_p0 = sext_ln126_1_fu_1662_p1;
  assign grp_fu_4473_p1 = sext_ln105_1_reg_4871;
  assign grp_fu_4481_p0 = sext_ln126_1_fu_1662_p1;
  assign grp_fu_4481_p1 = sext_ln100_1_reg_4854;
  assign grp_fu_4489_p0 = sext_ln126_1_fu_1662_p1;
  assign grp_fu_4489_p1 = sext_ln96_1_reg_4836;
  assign grp_fu_4497_p0 = sext_ln126_1_fu_1662_p1;
  assign grp_fu_4497_p1 = sext_ln93_1_reg_4818;
  assign Const_754 = (16'd61082 ^ working_key[1977:1962]);
  assign grp_fu_4555_p2 = Const_754;
  assign grp_fu_4564_p1 = sext_ln62_2_reg_5457;
  assign Const_755 = (16'd2394 ^ working_key[1993:1978]);
  assign grp_fu_4564_p2 = Const_755;
  assign grp_fu_4572_p0 = sext_ln62_2_reg_5457;
  assign Const_756 = (16'd48437 ^ working_key[2009:1994]);
  assign grp_fu_4572_p2 = Const_756;
  assign Const_757 = (4'd4 ^ working_key[2013:2010]);
  assign i_1_fu_2491_p2 = (working_key[2014] == 1'b1)? i_2_i_reg_939 + Const_757 : i_2_i_reg_939 * Const_757;
  assign Const_758 = (4'd3 ^ working_key[2018:2015]);
  assign i_2_fu_2503_p2 = (working_key[2019] == 1'b1)? i_3_i_reg_950 + Const_758 : i_3_i_reg_950 - Const_758;
  assign Const_759 = (4'd11 ^ working_key[2023:2020]);
  assign i_fu_2449_p2 = (working_key[2024] == 1'b1)? i_1_i_reg_928 << Const_759 : i_1_i_reg_928 + Const_759;
  assign Const_760 = (64'd7660633594411619668 ^ working_key[2088:2025]);
  assign Const_761 = (1'd1 ^ working_key[2090]);
  assign Const_762 = (1'd1 ^ working_key[2091]);
  assign icmp_ln118_1_fu_2107_p2 = ((((working_key[2089] == 1'b1)? L_ACF_q0 != Const_760 : L_ACF_q0 < Const_760) ^ working_key[2092]) == 1'b1)? Const_761 : Const_762;
  assign Const_763 = (32'd1387617588 ^ working_key[2124:2093]);
  assign Const_764 = (1'd0 ^ working_key[2126]);
  assign Const_765 = (1'd0 ^ working_key[2127]);
  assign icmp_ln118_fu_1151_p2 = ((((working_key[2125] == 1'b1)? a_assign_1_fu_1143_p3 != Const_763 : a_assign_1_fu_1143_p3 < Const_763) ^ working_key[2128]) == 1'b1)? Const_765 : Const_764;
  assign Const_766 = (8'd166 ^ working_key[2136:2129]);
  assign Const_767 = (1'd0 ^ working_key[2138]);
  assign Const_768 = (1'd1 ^ working_key[2139]);
  assign icmp_ln123_1_fu_1231_p2 = ((((working_key[2137] == 1'b1)? tmp_3_fu_1221_p4 == Const_766 : tmp_3_fu_1221_p4 != Const_766) ^ working_key[2140]) == 1'b1)? Const_768 : Const_767;
  assign Const_769 = (24'd5592235 ^ working_key[2164:2141]);
  assign Const_770 = (1'd1 ^ working_key[2166]);
  assign Const_771 = (1'd1 ^ working_key[2167]);
  assign icmp_ln123_2_fu_1286_p2 = ((((working_key[2165] == 1'b1)? tmp_4_fu_1276_p4 == Const_769 : tmp_4_fu_1276_p4 > Const_769) ^ working_key[2168]) == 1'b1)? Const_770 : Const_771;
  assign Const_772 = (16'd21825 ^ working_key[2184:2169]);
  assign Const_773 = (1'd1 ^ working_key[2186]);
  assign Const_774 = (1'd1 ^ working_key[2187]);
  assign icmp_ln123_3_fu_2203_p2 = ((((working_key[2185] == 1'b1)? tmp_17_fu_2193_p4 == Const_772 : tmp_17_fu_2193_p4 === Const_772) ^ working_key[2188]) == 1'b1)? Const_773 : Const_774;
  assign Const_775 = (8'd85 ^ working_key[2196:2189]);
  assign Const_776 = (1'd0 ^ working_key[2198]);
  assign Const_777 = (1'd1 ^ working_key[2199]);
  assign icmp_ln123_4_fu_2219_p2 = ((((working_key[2197] == 1'b1)? tmp_18_fu_2209_p4 > Const_775 : tmp_18_fu_2209_p4 == Const_775) ^ working_key[2200]) == 1'b1)? Const_776 : Const_777;
  assign Const_778 = (1'd0 ^ working_key[2201]);
  assign Const_779 = (1'd1 ^ working_key[2203]);
  assign Const_780 = (1'd1 ^ working_key[2204]);
  assign icmp_ln123_5_fu_2309_p2 = ((((working_key[2202] == 1'b1)? tmp_19_fu_2299_p4 != Const_778 : tmp_19_fu_2299_p4 === Const_778) ^ working_key[2205]) == 1'b1)? Const_779 : Const_780;
  assign Const_781 = (24'd10134701 ^ working_key[2229:2206]);
  assign Const_782 = (1'd0 ^ working_key[2231]);
  assign Const_783 = (1'd1 ^ working_key[2232]);
  assign icmp_ln123_6_fu_2337_p2 = ((((working_key[2230] == 1'b1)? tmp_20_fu_2327_p4 > Const_781 : tmp_20_fu_2327_p4 == Const_781) ^ working_key[2233]) == 1'b1)? Const_783 : Const_782;
  assign Const_784 = (16'd38314 ^ working_key[2249:2234]);
  assign Const_785 = (1'd1 ^ working_key[2251]);
  assign Const_786 = (1'd1 ^ working_key[2252]);
  assign icmp_ln123_fu_1215_p2 = ((((working_key[2250] == 1'b1)? tmp_2_fu_1205_p4 === Const_784 : tmp_2_fu_1205_p4 == Const_784) ^ working_key[2253]) == 1'b1)? Const_785 : Const_786;
  assign Const_787 = (8'd173 ^ working_key[2261:2254]);
  assign Const_788 = (1'd1 ^ working_key[2263]);
  assign Const_789 = (1'd1 ^ working_key[2264]);
  assign icmp_ln135_fu_1848_p2 = ((((working_key[2262] == 1'b1)? sp_0_rec_i_reg_894 == Const_787 : sp_0_rec_i_reg_894 < Const_787) ^ working_key[2265]) == 1'b1)? Const_789 : Const_788;
  assign Const_790 = (16'd42335 ^ working_key[2281:2266]);
  assign Const_791 = (1'd0 ^ working_key[2283]);
  assign Const_792 = (1'd0 ^ working_key[2284]);
  assign icmp_ln147_fu_2573_p2 = ((((working_key[2282] == 1'b1)? temp_24_reg_997 < Const_790 : temp_24_reg_997 == Const_790) ^ working_key[2285]) == 1'b1)? Const_792 : Const_791;
  assign Const_793 = (4'd10 ^ working_key[2289:2286]);
  assign Const_794 = (1'd0 ^ working_key[2291]);
  assign Const_795 = (1'd0 ^ working_key[2292]);
  assign icmp_ln150_fu_2589_p2 = ((((working_key[2290] == 1'b1)? k_0_i_i_reg_1026 < Const_793 : k_0_i_i_reg_1026 == Const_793) ^ working_key[2293]) == 1'b1)? Const_795 : Const_794;
  assign Const_796 = (1'd0 ^ working_key[2295]);
  assign Const_797 = (1'd0 ^ working_key[2296]);
  assign icmp_ln155_fu_2601_p2 = ((((working_key[2294] == 1'b1)? L_num_1_fu_2595_p2 > sext_ln139_reg_5396 : L_num_1_fu_2595_p2 < sext_ln139_reg_5396) ^ working_key[2297]) == 1'b1)? Const_797 : Const_796;
  assign Const_798 = (8'd0 ^ working_key[2305:2298]);
  assign Const_799 = (1'd0 ^ working_key[2307]);
  assign Const_800 = (1'd0 ^ working_key[2308]);
  assign icmp_ln158_fu_2083_p2 = ((((working_key[2306] == 1'b1)? p_0_rec_i_reg_917 != Const_798 : p_0_rec_i_reg_917 == Const_798) ^ working_key[2309]) == 1'b1)? Const_800 : Const_799;
  assign Const_801 = (64'd6534330141437012650 ^ working_key[2373:2310]);
  assign Const_802 = (1'd1 ^ working_key[2375]);
  assign Const_803 = (1'd0 ^ working_key[2376]);
  assign icmp_ln178_fu_2101_p2 = ((((working_key[2374] == 1'b1)? L_ACF_q0 == Const_801 : L_ACF_q0 > Const_801) ^ working_key[2377]) == 1'b1)? Const_803 : Const_802;
  assign Const_804 = (4'd12 ^ working_key[2381:2378]);
  assign Const_805 = (1'd1 ^ working_key[2383]);
  assign Const_806 = (1'd1 ^ working_key[2384]);
  assign icmp_ln180_fu_3008_p2 = ((((working_key[2382] == 1'b1)? p_0_rec_i1_reg_1071 == Const_804 : p_0_rec_i1_reg_1071 > Const_804) ^ working_key[2385]) == 1'b1)? Const_805 : Const_806;
  assign Const_807 = (4'd10 ^ working_key[2389:2386]);
  assign Const_808 = (1'd1 ^ working_key[2391]);
  assign Const_809 = (1'd1 ^ working_key[2392]);
  assign icmp_ln186_fu_2443_p2 = ((((working_key[2390] == 1'b1)? i_1_i_reg_928 == Const_807 : i_1_i_reg_928 != Const_807) ^ working_key[2393]) == 1'b1)? Const_809 : Const_808;
  assign Const_810 = (4'd7 ^ working_key[2397:2394]);
  assign Const_811 = (1'd1 ^ working_key[2399]);
  assign Const_812 = (1'd1 ^ working_key[2400]);
  assign icmp_ln192_fu_2480_p2 = ((((working_key[2398] == 1'b1)? i_2_i_reg_939 == Const_810 : i_2_i_reg_939 != Const_810) ^ working_key[2401]) == 1'b1)? Const_811 : Const_812;
  assign Const_813 = (4'd12 ^ working_key[2405:2402]);
  assign Const_814 = (1'd0 ^ working_key[2407]);
  assign Const_815 = (1'd0 ^ working_key[2408]);
  assign icmp_ln194_fu_2497_p2 = ((((working_key[2406] == 1'b1)? i_3_i_reg_950 != Const_813 : i_3_i_reg_950 == Const_813) ^ working_key[2409]) == 1'b1)? Const_815 : Const_814;
  assign icmp_ln204_fu_2555_p0 = P_q0;
  assign Const_816 = (1'd0 ^ working_key[2411]);
  assign Const_817 = (1'd0 ^ working_key[2412]);
  assign icmp_ln204_fu_2555_p2 = ((((working_key[2410] == 1'b1)? icmp_ln204_fu_2555_p0 == temp_24_reg_997 : icmp_ln204_fu_2555_p0 < temp_24_reg_997) ^ working_key[2413]) == 1'b1)? Const_817 : Const_816;
  assign Const_818 = (1'd0 ^ working_key[2415]);
  assign Const_819 = (1'd0 ^ working_key[2416]);
  assign icmp_ln206_fu_2677_p2 = ((((working_key[2414] == 1'b1)? p_2_rec_i_reg_1049 > indvars_iv142_reg_961 : p_2_rec_i_reg_1049 == indvars_iv142_reg_961) ^ working_key[2417]) == 1'b1)? Const_819 : Const_818;
  assign Const_820 = (16'd41130 ^ working_key[2433:2418]);
  assign Const_821 = (1'd0 ^ working_key[2435]);
  assign Const_822 = (1'd0 ^ working_key[2436]);
  assign icmp_ln213_fu_2637_p2 = ((((working_key[2434] == 1'b1)? temp_3_reg_5366 == Const_820 : temp_3_reg_5366 > Const_820) ^ working_key[2437]) == 1'b1)? Const_822 : Const_821;
  assign Const_823 = (32'd2907908770 ^ working_key[2469:2438]);
  assign Const_824 = (1'd1 ^ working_key[2471]);
  assign Const_825 = (1'd1 ^ working_key[2472]);
  assign icmp_ln215_fu_2657_p2 = ((((working_key[2470] == 1'b1)? i_3_reg_973 != Const_823 : i_3_reg_973 == Const_823) ^ working_key[2473]) == 1'b1)? Const_824 : Const_825;
  assign Const_826 = (1'd0 ^ working_key[2475]);
  assign Const_827 = (1'd0 ^ working_key[2476]);
  assign icmp_ln223_fu_2788_p2 = ((((working_key[2474] == 1'b1)? m_0_i_reg_1060 < sub_ln223_reg_5468 : m_0_i_reg_1060 > sub_ln223_reg_5468) ^ working_key[2477]) == 1'b1)? Const_827 : Const_826;
  assign Const_828 = (4'd2 ^ working_key[2481:2478]);
  assign Const_829 = (1'd1 ^ working_key[2483]);
  assign Const_830 = (1'd0 ^ working_key[2484]);
  assign icmp_ln253_fu_3025_p2 = ((((working_key[2482] == 1'b1)? p_0_rec_i16_reg_1082 == Const_828 : p_0_rec_i16_reg_1082 < Const_828) ^ working_key[2485]) == 1'b1)? Const_830 : Const_829;
  assign Const_831 = (16'd3272 ^ working_key[2501:2486]);
  assign Const_832 = (1'd1 ^ working_key[2503]);
  assign Const_833 = (1'd0 ^ working_key[2504]);
  assign icmp_ln259_fu_3073_p2 = ((((working_key[2502] == 1'b1)? temp_fu_3065_p3 < Const_831 : temp_fu_3065_p3 === Const_831) ^ working_key[2505]) == 1'b1)? Const_833 : Const_832;
  assign Const_834 = (16'd43726 ^ working_key[2521:2506]);
  assign Const_835 = (1'd0 ^ working_key[2523]);
  assign Const_836 = (1'd1 ^ working_key[2524]);
  assign icmp_ln263_fu_3093_p2 = ((((working_key[2522] == 1'b1)? temp_fu_3065_p3 < Const_834 : temp_fu_3065_p3 > Const_834) ^ working_key[2525]) == 1'b1)? Const_836 : Const_835;
  assign Const_837 = (7'd53 ^ working_key[2532:2526]);
  assign Const_838 = (1'd1 ^ working_key[2534]);
  assign Const_839 = (1'd1 ^ working_key[2535]);
  assign icmp_ln304_1_fu_3628_p2 = ((((working_key[2533] == 1'b1)? select_ln40_6_fu_3602_p3 === Const_837 : select_ln40_6_fu_3602_p3 < Const_837) ^ working_key[2536]) == 1'b1)? Const_838 : Const_839;
  assign Const_840 = (2'd0 ^ working_key[2538:2537]);
  assign Const_841 = (1'd1 ^ working_key[2540]);
  assign Const_842 = (1'd1 ^ working_key[2541]);
  assign icmp_ln304_fu_3622_p2 = ((((working_key[2539] == 1'b1)? tmp_26_fu_3612_p4 == Const_840 : tmp_26_fu_3612_p4 != Const_840) ^ working_key[2542]) == 1'b1)? Const_841 : Const_842;
  assign Const_843 = (7'd53 ^ working_key[2549:2543]);
  assign Const_844 = (1'd0 ^ working_key[2551]);
  assign Const_845 = (1'd0 ^ working_key[2552]);
  assign icmp_ln305_1_fu_3693_p2 = ((((working_key[2550] == 1'b1)? select_ln40_7_fu_3667_p3 == Const_843 : select_ln40_7_fu_3667_p3 < Const_843) ^ working_key[2553]) == 1'b1)? Const_845 : Const_844;
  assign Const_846 = (2'd1 ^ working_key[2555:2554]);
  assign Const_847 = (1'd1 ^ working_key[2557]);
  assign Const_848 = (1'd0 ^ working_key[2558]);
  assign icmp_ln305_fu_3687_p2 = ((((working_key[2556] == 1'b1)? tmp_28_fu_3677_p4 < Const_846 : tmp_28_fu_3677_p4 == Const_846) ^ working_key[2559]) == 1'b1)? Const_848 : Const_847;
  assign Const_849 = (7'd90 ^ working_key[2566:2560]);
  assign Const_850 = (1'd1 ^ working_key[2568]);
  assign Const_851 = (1'd1 ^ working_key[2569]);
  assign icmp_ln306_1_fu_3864_p2 = ((((working_key[2567] == 1'b1)? select_ln40_9_fu_3838_p3 < Const_849 : select_ln40_9_fu_3838_p3 > Const_849) ^ working_key[2570]) == 1'b1)? Const_850 : Const_851;
  assign Const_852 = (3'd5 ^ working_key[2573:2571]);
  assign Const_853 = (1'd0 ^ working_key[2575]);
  assign Const_854 = (1'd0 ^ working_key[2576]);
  assign icmp_ln306_fu_3858_p2 = ((((working_key[2574] == 1'b1)? tmp_31_fu_3848_p4 === Const_852 : tmp_31_fu_3848_p4 > Const_852) ^ working_key[2577]) == 1'b1)? Const_854 : Const_853;
  assign Const_855 = (7'd66 ^ working_key[2584:2578]);
  assign Const_856 = (1'd0 ^ working_key[2586]);
  assign Const_857 = (1'd0 ^ working_key[2587]);
  assign icmp_ln307_1_fu_3929_p2 = ((((working_key[2585] == 1'b1)? select_ln40_10_fu_3903_p3 === Const_855 : select_ln40_10_fu_3903_p3 < Const_855) ^ working_key[2588]) == 1'b1)? Const_857 : Const_856;
  assign Const_858 = (3'd5 ^ working_key[2591:2589]);
  assign Const_859 = (1'd0 ^ working_key[2593]);
  assign Const_860 = (1'd0 ^ working_key[2594]);
  assign icmp_ln307_fu_3923_p2 = ((((working_key[2592] == 1'b1)? tmp_32_fu_3913_p4 === Const_858 : tmp_32_fu_3913_p4 > Const_858) ^ working_key[2595]) == 1'b1)? Const_859 : Const_860;
  assign Const_861 = (7'd81 ^ working_key[2602:2596]);
  assign Const_862 = (1'd1 ^ working_key[2604]);
  assign Const_863 = (1'd1 ^ working_key[2605]);
  assign icmp_ln309_1_fu_4054_p2 = ((((working_key[2603] == 1'b1)? select_ln40_12_fu_4028_p3 < Const_861 : select_ln40_12_fu_4028_p3 === Const_861) ^ working_key[2606]) == 1'b1)? Const_863 : Const_862;
  assign Const_864 = (4'd4 ^ working_key[2610:2607]);
  assign Const_865 = (1'd0 ^ working_key[2612]);
  assign Const_866 = (1'd1 ^ working_key[2613]);
  assign icmp_ln309_fu_4048_p2 = ((((working_key[2611] == 1'b1)? tmp_35_fu_4038_p4 > Const_864 : tmp_35_fu_4038_p4 < Const_864) ^ working_key[2614]) == 1'b1)? Const_865 : Const_866;
  assign Const_867 = (7'd45 ^ working_key[2621:2615]);
  assign Const_868 = (1'd1 ^ working_key[2623]);
  assign Const_869 = (1'd1 ^ working_key[2624]);
  assign icmp_ln310_1_fu_4119_p2 = ((((working_key[2622] == 1'b1)? select_ln40_13_fu_4093_p3 < Const_867 : select_ln40_13_fu_4093_p3 > Const_867) ^ working_key[2625]) == 1'b1)? Const_868 : Const_869;
  assign Const_870 = (4'd9 ^ working_key[2629:2626]);
  assign Const_871 = (1'd1 ^ working_key[2631]);
  assign Const_872 = (1'd1 ^ working_key[2632]);
  assign icmp_ln310_fu_4113_p2 = ((((working_key[2630] == 1'b1)? tmp_36_fu_4103_p4 < Const_870 : tmp_36_fu_4103_p4 > Const_870) ^ working_key[2633]) == 1'b1)? Const_871 : Const_872;
  assign Const_873 = (7'd73 ^ working_key[2640:2634]);
  assign Const_874 = (1'd0 ^ working_key[2642]);
  assign Const_875 = (1'd0 ^ working_key[2643]);
  assign icmp_ln311_1_fu_4184_p2 = ((((working_key[2641] == 1'b1)? select_ln40_14_fu_4158_p3 === Const_873 : select_ln40_14_fu_4158_p3 < Const_873) ^ working_key[2644]) == 1'b1)? Const_875 : Const_874;
  assign Const_876 = (5'd31 ^ working_key[2649:2645]);
  assign Const_877 = (1'd1 ^ working_key[2651]);
  assign Const_878 = (1'd1 ^ working_key[2652]);
  assign icmp_ln311_fu_4178_p2 = ((((working_key[2650] == 1'b1)? tmp_37_fu_4168_p4 > Const_876 : tmp_37_fu_4168_p4 != Const_876) ^ working_key[2653]) == 1'b1)? Const_877 : Const_878;
  assign Const_879 = (7'd89 ^ working_key[2660:2654]);
  assign Const_880 = (1'd1 ^ working_key[2662]);
  assign Const_881 = (1'd1 ^ working_key[2663]);
  assign icmp_ln312_1_fu_4249_p2 = ((((working_key[2661] == 1'b1)? select_ln40_15_fu_4223_p3 < Const_879 : select_ln40_15_fu_4223_p3 === Const_879) ^ working_key[2664]) == 1'b1)? Const_880 : Const_881;
  assign Const_882 = (5'd21 ^ working_key[2669:2665]);
  assign Const_883 = (1'd0 ^ working_key[2671]);
  assign Const_884 = (1'd0 ^ working_key[2672]);
  assign icmp_ln312_fu_4243_p2 = ((((working_key[2670] == 1'b1)? tmp_38_fu_4233_p4 === Const_882 : tmp_38_fu_4233_p4 > Const_882) ^ working_key[2673]) == 1'b1)? Const_884 : Const_883;
  assign Const_885 = (2'd3 ^ working_key[2675:2674]);
  assign Const_886 = (1'd0 ^ working_key[2677]);
  assign Const_887 = (1'd0 ^ working_key[2678]);
  assign icmp_ln40_10_fu_3423_p2 = ((((working_key[2676] == 1'b1)? tmp_30_fu_3413_p4 > Const_885 : tmp_30_fu_3413_p4 == Const_885) ^ working_key[2679]) == 1'b1)? Const_886 : Const_887;
  assign Const_888 = (2'd1 ^ working_key[2681:2680]);
  assign Const_889 = (1'd0 ^ working_key[2683]);
  assign Const_890 = (1'd0 ^ working_key[2684]);
  assign icmp_ln40_11_fu_3751_p2 = ((((working_key[2682] == 1'b1)? tmp_33_fu_3741_p4 > Const_888 : tmp_33_fu_3741_p4 == Const_888) ^ working_key[2685]) == 1'b1)? Const_890 : Const_889;
  assign Const_891 = (2'd3 ^ working_key[2687:2686]);
  assign Const_892 = (1'd0 ^ working_key[2689]);
  assign Const_893 = (1'd0 ^ working_key[2690]);
  assign icmp_ln40_12_fu_3790_p2 = ((((working_key[2688] == 1'b1)? tmp_34_fu_3780_p4 > Const_891 : tmp_34_fu_3780_p4 == Const_891) ^ working_key[2691]) == 1'b1)? Const_893 : Const_892;
  assign Const_894 = (17'd84650 ^ working_key[2708:2692]);
  assign Const_895 = (1'd0 ^ working_key[2710]);
  assign Const_896 = (1'd0 ^ working_key[2711]);
  assign icmp_ln40_13_fu_3580_p2 = ((((working_key[2709] == 1'b1)? sum_10_fu_3574_p2 != Const_894 : sum_10_fu_3574_p2 < Const_894) ^ working_key[2712]) == 1'b1)? Const_896 : Const_895;
  assign Const_897 = (17'd51546 ^ working_key[2729:2713]);
  assign Const_898 = (1'd0 ^ working_key[2731]);
  assign Const_899 = (1'd0 ^ working_key[2732]);
  assign icmp_ln40_14_fu_3977_p2 = ((((working_key[2730] == 1'b1)? sum_11_fu_3971_p2 != Const_897 : sum_11_fu_3971_p2 < Const_897) ^ working_key[2733]) == 1'b1)? Const_899 : Const_898;
  assign Const_900 = (17'd10985 ^ working_key[2750:2734]);
  assign Const_901 = (1'd0 ^ working_key[2752]);
  assign Const_902 = (1'd0 ^ working_key[2753]);
  assign icmp_ln40_15_fu_4007_p2 = ((((working_key[2751] == 1'b1)? sum_12_fu_4001_p2 > Const_900 : sum_12_fu_4001_p2 < Const_900) ^ working_key[2754]) == 1'b1)? Const_902 : Const_901;
  assign Const_903 = (2'd1 ^ working_key[2756:2755]);
  assign Const_904 = (1'd1 ^ working_key[2758]);
  assign Const_905 = (1'd0 ^ working_key[2759]);
  assign icmp_ln40_1_fu_2748_p2 = ((((working_key[2757] == 1'b1)? tmp_22_fu_2738_p4 == Const_903 : tmp_22_fu_2738_p4 === Const_903) ^ working_key[2760]) == 1'b1)? Const_905 : Const_904;
  assign Const_906 = (17'd31338 ^ working_key[2777:2761]);
  assign Const_907 = (1'd1 ^ working_key[2779]);
  assign Const_908 = (1'd1 ^ working_key[2780]);
  assign icmp_ln40_2_fu_2895_p2 = ((((working_key[2778] == 1'b1)? sum_1_fu_2889_p2 < Const_906 : sum_1_fu_2889_p2 === Const_906) ^ working_key[2781]) == 1'b1)? Const_907 : Const_908;
  assign Const_909 = (2'd0 ^ working_key[2783:2782]);
  assign Const_910 = (1'd1 ^ working_key[2785]);
  assign Const_911 = (1'd0 ^ working_key[2786]);
  assign icmp_ln40_3_fu_2911_p2 = ((((working_key[2784] == 1'b1)? tmp_23_fu_2901_p4 == Const_909 : tmp_23_fu_2901_p4 != Const_909) ^ working_key[2787]) == 1'b1)? Const_911 : Const_910;
  assign Const_912 = (17'd76458 ^ working_key[2804:2788]);
  assign Const_913 = (1'd1 ^ working_key[2806]);
  assign Const_914 = (1'd0 ^ working_key[2807]);
  assign icmp_ln40_4_fu_2954_p2 = ((((working_key[2805] == 1'b1)? sum_2_fu_2948_p2 < Const_912 : sum_2_fu_2948_p2 != Const_912) ^ working_key[2808]) == 1'b1)? Const_913 : Const_914;
  assign Const_915 = (2'd1 ^ working_key[2810:2809]);
  assign Const_916 = (1'd1 ^ working_key[2812]);
  assign Const_917 = (1'd1 ^ working_key[2813]);
  assign icmp_ln40_5_fu_2970_p2 = ((((working_key[2811] == 1'b1)? tmp_24_fu_2960_p4 == Const_915 : tmp_24_fu_2960_p4 < Const_915) ^ working_key[2814]) == 1'b1)? Const_916 : Const_917;
  assign Const_918 = (2'd0 ^ working_key[2816:2815]);
  assign Const_919 = (1'd1 ^ working_key[2818]);
  assign Const_920 = (1'd1 ^ working_key[2819]);
  assign icmp_ln40_6_fu_3219_p2 = ((((working_key[2817] == 1'b1)? tmp_25_fu_3209_p4 == Const_918 : tmp_25_fu_3209_p4 > Const_918) ^ working_key[2820]) == 1'b1)? Const_919 : Const_920;
  assign Const_921 = (2'd0 ^ working_key[2822:2821]);
  assign Const_922 = (1'd1 ^ working_key[2824]);
  assign Const_923 = (1'd1 ^ working_key[2825]);
  assign icmp_ln40_7_fu_3301_p2 = ((((working_key[2823] == 1'b1)? tmp_27_fu_3291_p4 == Const_921 : tmp_27_fu_3291_p4 != Const_921) ^ working_key[2826]) == 1'b1)? Const_922 : Const_923;
  assign Const_924 = (17'd81301 ^ working_key[2843:2827]);
  assign Const_925 = (1'd0 ^ working_key[2845]);
  assign Const_926 = (1'd0 ^ working_key[2846]);
  assign icmp_ln40_8_fu_3495_p2 = ((((working_key[2844] == 1'b1)? sum_7_fu_3489_p2 < Const_924 : sum_7_fu_3489_p2 == Const_924) ^ working_key[2847]) == 1'b1)? Const_926 : Const_925;
  assign Const_927 = (2'd3 ^ working_key[2849:2848]);
  assign Const_928 = (1'd1 ^ working_key[2851]);
  assign Const_929 = (1'd1 ^ working_key[2852]);
  assign icmp_ln40_9_fu_3383_p2 = ((((working_key[2850] == 1'b1)? tmp_29_fu_3373_p4 === Const_927 : tmp_29_fu_3373_p4 == Const_927) ^ working_key[2853]) == 1'b1)? Const_928 : Const_929;
  assign Const_930 = (17'd92586 ^ working_key[2870:2854]);
  assign Const_931 = (1'd1 ^ working_key[2872]);
  assign Const_932 = (1'd1 ^ working_key[2873]);
  assign icmp_ln40_fu_2732_p2 = ((((working_key[2871] == 1'b1)? sum_fu_2727_p2 < Const_930 : sum_fu_2727_p2 > Const_930) ^ working_key[2874]) == 1'b1)? Const_931 : Const_932;
  assign Const_933 = (16'd9389 ^ working_key[2890:2875]);
  assign Const_934 = (1'd0 ^ working_key[2892]);
  assign Const_935 = (1'd0 ^ working_key[2893]);
  assign icmp_ln58_1_fu_2689_p2 = ((((working_key[2891] == 1'b1)? select_ln213_reg_5434 < Const_933 : select_ln213_reg_5434 == Const_933) ^ working_key[2894]) == 1'b1)? Const_935 : Const_934;
  assign icmp_ln58_3_fu_2821_p0 = K_q0;
  assign Const_936 = (16'd12265 ^ working_key[2910:2895]);
  assign Const_937 = (1'd0 ^ working_key[2912]);
  assign Const_938 = (1'd0 ^ working_key[2913]);
  assign icmp_ln58_3_fu_2821_p2 = ((((working_key[2911] == 1'b1)? icmp_ln58_3_fu_2821_p0 != Const_936 : icmp_ln58_3_fu_2821_p0 == Const_936) ^ working_key[2914]) == 1'b1)? Const_937 : Const_938;
  assign Const_939 = (8'd245 ^ working_key[2922:2915]);
  assign Const_940 = (1'd1 ^ working_key[2924]);
  assign Const_941 = (1'd1 ^ working_key[2925]);
  assign icmp_ln58_fu_1126_p2 = ((((working_key[2923] == 1'b1)? k_0_i_reg_851 == Const_939 : k_0_i_reg_851 != Const_939) ^ working_key[2926]) == 1'b1)? Const_940 : Const_941;
  assign Const_942 = (1'd1 ^ working_key[2928]);
  assign Const_943 = (1'd1 ^ working_key[2929]);
  assign icmp_ln61_fu_1328_p2 = ((((working_key[2927] == 1'b1)? smax_fu_1320_p3 > smax_0_i_reg_839 : smax_fu_1320_p3 != smax_0_i_reg_839) ^ working_key[2930]) == 1'b1)? Const_942 : Const_943;
  assign Const_944 = (16'd21765 ^ working_key[2946:2931]);
  assign Const_945 = (1'd1 ^ working_key[2948]);
  assign Const_946 = (1'd1 ^ working_key[2949]);
  assign icmp_ln67_fu_1342_p2 = ((((working_key[2947] == 1'b1)? smax_0_i_reg_839 == Const_944 : smax_0_i_reg_839 < Const_944) ^ working_key[2950]) == 1'b1)? Const_945 : Const_946;
  assign Const_947 = (16'd6485 ^ working_key[2966:2951]);
  assign Const_948 = (1'd0 ^ working_key[2968]);
  assign Const_949 = (1'd0 ^ working_key[2969]);
  assign icmp_ln72_1_fu_1300_p2 = ((((working_key[2967] == 1'b1)? s_q0 != Const_947 : s_q0 == Const_947) ^ working_key[2970]) == 1'b1)? Const_949 : Const_948;
  assign Const_950 = (6'd19 ^ working_key[2976:2971]);
  assign Const_951 = (1'd1 ^ working_key[2978]);
  assign Const_952 = (1'd0 ^ working_key[2979]);
  assign icmp_ln72_2_fu_1489_p2 = ((((working_key[2977] == 1'b1)? n_fu_1471_p3 < Const_950 : n_fu_1471_p3 > Const_950) ^ working_key[2980]) == 1'b1)? Const_952 : Const_951;
  assign Const_953 = (16'd21332 ^ working_key[2996:2981]);
  assign Const_954 = (1'd1 ^ working_key[2998]);
  assign Const_955 = (1'd1 ^ working_key[2999]);
  assign icmp_ln72_4_fu_3045_p2 = ((((working_key[2997] == 1'b1)? LARc_q0 == Const_953 : LARc_q0 === Const_953) ^ working_key[3000]) == 1'b1)? Const_954 : Const_955;
  assign Const_956 = (6'd53 ^ working_key[3006:3001]);
  assign Const_957 = (1'd0 ^ working_key[3008]);
  assign Const_958 = (1'd0 ^ working_key[3009]);
  assign icmp_ln72_fu_1483_p2 = ((((working_key[3007] == 1'b1)? n_fu_1471_p3 === Const_956 : n_fu_1471_p3 > Const_956) ^ working_key[3010]) == 1'b1)? Const_958 : Const_957;
  assign Const_959 = (8'd4 ^ working_key[3018:3011]);
  assign Const_960 = (1'd0 ^ working_key[3020]);
  assign Const_961 = (1'd0 ^ working_key[3021]);
  assign icmp_ln75_fu_1524_p2 = ((((working_key[3019] == 1'b1)? k_1_i_reg_862 != Const_959 : k_1_i_reg_862 == Const_959) ^ working_key[3022]) == 1'b1)? Const_961 : Const_960;
  assign Const_962 = (8'd232 ^ working_key[3030:3023]);
  assign k_1_fu_1530_p2 = (working_key[3031] == 1'b1)? k_1_i_reg_862 + Const_962 : k_1_i_reg_862 << Const_962;
  assign Const_963 = (5'd8 ^ working_key[3036:3032]);
  assign k_2_fu_1571_p2 = (working_key[3037] == 1'b1)? k_2_i_reg_873 << Const_963 : k_2_i_reg_873 + Const_963;
  assign Const_964 = (5'd26 ^ working_key[3042:3038]);
  assign k_3_fu_2065_p2 = (working_key[3043] == 1'b1)? Const_964 + k_3_i_reg_906 : Const_964 - k_3_i_reg_906;
  assign Const_965 = (8'd171 ^ working_key[3051:3044]);
  assign k_fu_1132_p2 = (working_key[3052] == 1'b1)? k_0_i_reg_851 << Const_965 : k_0_i_reg_851 + Const_965;
  assign Const_966 = (15'd341 ^ working_key[3067:3053]);
  assign lshr_ln76_fu_1514_p2 = (working_key[3068] == 1'b1)? Const_966 << zext_ln76_fu_1510_p1 : Const_966 >> zext_ln76_fu_1510_p1;
  assign Const_967 = (32'd2858767700 ^ working_key[3100:3069]);
  assign m_fu_2798_p2 = (working_key[3101] == 1'b1)? m_0_i_reg_1060 + Const_967 : m_0_i_reg_1060 << Const_967;
  assign mul_ln100_fu_4314_p0 = sext_ln100_1_fu_1596_p1;
  assign mul_ln100_fu_4314_p1 = sext_ln100_1_fu_1596_p1;
  assign mul_ln103_fu_4320_p0 = sext_ln100_1_fu_1596_p1;
  assign mul_ln103_fu_4320_p1 = sext_ln91_fu_1577_p1;
  assign mul_ln107_fu_4326_p0 = sext_ln105_1_fu_1599_p1;
  assign mul_ln107_fu_4326_p1 = sext_ln96_1_fu_1590_p1;
  assign mul_ln109_fu_4422_p0 = sext_ln105_1_reg_4871;
  assign mul_ln109_fu_4422_p1 = sext_ln91_reg_4810;
  assign mul_ln111_fu_4426_p0 = sext_ln111_1_reg_4896;
  assign mul_ln111_fu_4426_p1 = sext_ln111_1_reg_4896;
  assign mul_ln116_fu_4332_p1 = sext_ln91_fu_1577_p1;
  assign mul_ln118_fu_4338_p0 = sext_ln118_1_fu_1612_p1;
  assign mul_ln118_fu_4338_p1 = sext_ln118_1_fu_1612_p1;
  assign mul_ln120_fu_4344_p0 = sext_ln118_1_fu_1612_p1;
  assign mul_ln120_fu_4344_p1 = sext_ln105_1_fu_1599_p1;
  assign mul_ln121_fu_4350_p0 = sext_ln118_1_fu_1612_p1;
  assign mul_ln121_fu_4350_p1 = sext_ln100_1_fu_1596_p1;
  assign mul_ln122_fu_4356_p0 = sext_ln118_1_fu_1612_p1;
  assign mul_ln122_fu_4356_p1 = sext_ln96_1_fu_1590_p1;
  assign mul_ln123_fu_4362_p0 = sext_ln118_1_fu_1612_p1;
  assign mul_ln123_fu_4362_p1 = sext_ln93_1_fu_1584_p1;
  assign mul_ln124_fu_4368_p0 = sext_ln118_1_fu_1612_p1;
  assign mul_ln124_fu_4368_p1 = sext_ln91_fu_1577_p1;
  assign mul_ln133_fu_4504_p0 = sext_ln126_1_fu_1662_p1;
  assign mul_ln133_fu_4504_p1 = sext_ln91_reg_4810;
  assign mul_ln140_fu_4521_p0 = sext_ln140_reg_5089;
  assign mul_ln140_fu_4521_p1 = sext_ln140_reg_5089;
  assign mul_ln141_fu_4509_p1 = sext_ln140_fu_1882_p1;
  assign mul_ln142_fu_4515_p1 = sext_ln140_fu_1882_p1;
  assign mul_ln143_fu_4525_p1 = sext_ln140_reg_5089;
  assign mul_ln144_fu_4530_p1 = sext_ln140_reg_5089;
  assign mul_ln145_fu_4535_p1 = sext_ln140_reg_5089;
  assign mul_ln146_fu_4540_p1 = sext_ln140_reg_5089;
  assign mul_ln147_fu_4545_p1 = sext_ln140_reg_5089;
  assign mul_ln148_fu_4550_p1 = sext_ln140_reg_5089;
  assign Const_968 = (15'd2844 ^ working_key[3116:3102]);
  assign mul_ln50_1_fu_4587_p1 = Const_968;
  assign Const_969 = (15'd30367 ^ working_key[3131:3117]);
  assign mul_ln50_2_fu_4594_p1 = Const_969;
  assign Const_970 = (15'd25818 ^ working_key[3146:3132]);
  assign mul_ln50_fu_4580_p1 = Const_970;
  assign mul_ln93_fu_4296_p0 = sext_ln93_1_fu_1584_p1;
  assign mul_ln93_fu_4296_p1 = sext_ln93_1_fu_1584_p1;
  assign mul_ln94_fu_4302_p0 = sext_ln93_1_fu_1584_p1;
  assign mul_ln94_fu_4302_p1 = sext_ln91_fu_1577_p1;
  assign mul_ln98_fu_4308_p0 = sext_ln96_1_fu_1590_p1;
  assign mul_ln98_fu_4308_p1 = sext_ln91_fu_1577_p1;
  assign Const_971 = (32'd1428881051 ^ working_key[3178:3147]);
  assign n_1_fu_2809_p2 = (working_key[3179] == 1'b1)? i_3_reg_973 + Const_971 : i_3_reg_973 << Const_971;
  assign Const_972 = (1'd1 ^ working_key[3180]);
  assign n_fu_1471_p3 = ((((working_key[3181] == 1'b1)? or_ln67_fu_1466_p2[0:0] === Const_972 : or_ln67_fu_1466_p2[0:0] > Const_972) ^ working_key[3182]) == 1'b1)? select_ln67_fu_1458_p3 : sub_ln70_fu_1452_p2;
  assign newSel112_cast_fu_1440_p1 = newSel112_fu_1432_p3;
  assign Const_973 = (1'd0 ^ working_key[3183]);
  assign newSel112_fu_1432_p3 = ((((working_key[3184] == 1'b1)? sel_tmp24_fu_1388_p2[0:0] != Const_973 : sel_tmp24_fu_1388_p2[0:0] === Const_973) ^ working_key[3185]) == 1'b1)? sext_ln123_fu_1368_p1 : zext_ln123_2_fu_1358_p1;
  assign Const_974 = (1'd1 ^ working_key[3186]);
  assign newSel114_fu_1444_p3 = ((((working_key[3187] == 1'b1)? or_cond_fu_1426_p2[0:0] === Const_974 : or_cond_fu_1426_p2[0:0] == Const_974) ^ working_key[3188]) == 1'b1)? newSel_cast_fu_1422_p1 : newSel112_cast_fu_1440_p1;
  assign newSel_cast_fu_1422_p1 = newSel_fu_1416_p2;
  assign newSel_fu_1416_p2 = (working_key[3189] == 1'b1)? zext_ln123_fu_1348_p1 + newSel_v_fu_1408_p3 : zext_ln123_fu_1348_p1 * newSel_v_fu_1408_p3;
  assign Const_975 = (1'd1 ^ working_key[3190]);
  assign Const_976 = (5'd31 ^ working_key[3196:3192]);
  assign Const_977 = (5'd26 ^ working_key[3201:3197]);
  assign newSel_v_fu_1408_p3 = ((((working_key[3191] == 1'b1)? sel_tmp37_fu_1403_p2[0:0] > Const_975 : sel_tmp37_fu_1403_p2[0:0] === Const_975) ^ working_key[3202]) == 1'b1)? Const_976 : Const_977;
  assign or_cond_fu_1426_p2 = (working_key[3203] == 1'b1)? sel_tmp37_fu_1403_p2 | sel_tmp31_fu_1398_p2 : sel_tmp37_fu_1403_p2 ^ sel_tmp31_fu_1398_p2;
  assign or_ln118_1_fu_2355_p2 = (working_key[3204] == 1'b1)? sel_tmp57_fu_2321_p2 >> sel_tmp50_fu_2293_p2 : sel_tmp57_fu_2321_p2 | sel_tmp50_fu_2293_p2;
  assign or_ln118_2_fu_2361_p2 = (working_key[3205] == 1'b1)? or_ln118_fu_2349_p2 | or_ln118_1_fu_2355_p2 : or_ln118_fu_2349_p2 << or_ln118_1_fu_2355_p2;
  assign or_ln118_fu_2349_p2 = (working_key[3206] == 1'b1)? sel_tmp63_fu_2343_p2 << icmp_ln118_1_fu_2107_p2 : sel_tmp63_fu_2343_p2 | icmp_ln118_1_fu_2107_p2;
  assign or_ln304_fu_3648_p2 = (working_key[3207] == 1'b1)? icmp_ln304_fu_3622_p2 | icmp_ln304_1_fu_3628_p2 : icmp_ln304_fu_3622_p2 << icmp_ln304_1_fu_3628_p2;
  assign or_ln305_fu_3713_p2 = (working_key[3208] == 1'b1)? icmp_ln305_fu_3687_p2 ^ icmp_ln305_1_fu_3693_p2 : icmp_ln305_fu_3687_p2 | icmp_ln305_1_fu_3693_p2;
  assign or_ln306_fu_3884_p2 = (working_key[3209] == 1'b1)? icmp_ln306_fu_3858_p2 | icmp_ln306_1_fu_3864_p2 : icmp_ln306_fu_3858_p2 << icmp_ln306_1_fu_3864_p2;
  assign or_ln307_fu_3949_p2 = (working_key[3210] == 1'b1)? icmp_ln307_fu_3923_p2 & icmp_ln307_1_fu_3929_p2 : icmp_ln307_fu_3923_p2 | icmp_ln307_1_fu_3929_p2;
  assign or_ln309_fu_4074_p2 = (working_key[3211] == 1'b1)? icmp_ln309_fu_4048_p2 | icmp_ln309_1_fu_4054_p2 : icmp_ln309_fu_4048_p2 << icmp_ln309_1_fu_4054_p2;
  assign or_ln310_fu_4139_p2 = (working_key[3212] == 1'b1)? icmp_ln310_fu_4113_p2 & icmp_ln310_1_fu_4119_p2 : icmp_ln310_fu_4113_p2 | icmp_ln310_1_fu_4119_p2;
  assign or_ln311_fu_4204_p2 = (working_key[3213] == 1'b1)? icmp_ln311_fu_4178_p2 | icmp_ln311_1_fu_4184_p2 : icmp_ln311_fu_4178_p2 & icmp_ln311_1_fu_4184_p2;
  assign or_ln312_fu_4269_p2 = (working_key[3214] == 1'b1)? icmp_ln312_fu_4243_p2 >> icmp_ln312_1_fu_4249_p2 : icmp_ln312_fu_4243_p2 | icmp_ln312_1_fu_4249_p2;
  assign or_ln40_1_fu_2930_p2 = (working_key[3215] == 1'b1)? icmp_ln40_3_fu_2911_p2 | icmp_ln40_2_fu_2895_p2 : icmp_ln40_3_fu_2911_p2 >> icmp_ln40_2_fu_2895_p2;
  assign or_ln40_2_fu_2988_p2 = (working_key[3216] == 1'b1)? icmp_ln40_5_fu_2970_p2 & icmp_ln40_4_fu_2954_p2 : icmp_ln40_5_fu_2970_p2 | icmp_ln40_4_fu_2954_p2;
  assign or_ln40_fu_2768_p2 = (working_key[3217] == 1'b1)? icmp_ln40_fu_2732_p2 << icmp_ln40_1_fu_2748_p2 : icmp_ln40_fu_2732_p2 | icmp_ln40_1_fu_2748_p2;
  assign or_ln67_fu_1466_p2 = (working_key[3218] == 1'b1)? icmp_ln67_fu_1342_p2 | icmp_ln118_reg_4631 : icmp_ln67_fu_1342_p2 >> icmp_ln118_reg_4631;
  assign p_0_rec_i16_cast_fu_3020_p1 = p_0_rec_i16_reg_1082;
  assign p_0_rec_i1_cast_fu_3003_p1 = p_0_rec_i1_reg_1071;
  assign p_0_rec_i_cast_fu_2078_p1 = p_0_rec_i_reg_917;
  assign s_d0 = trunc_ln2_reg_4714;
  assign s_d1 = (working_key[3219] == 1'b1)? s_q1 << sext_ln67_reg_4678 : s_q1 >> sext_ln67_reg_4678;
  assign sel_tmp24_fu_1388_p2 = (working_key[3220] == 1'b1)? tmp_fu_1382_p2 | icmp_ln123_1_reg_4648 : tmp_fu_1382_p2 & icmp_ln123_1_reg_4648;
  assign sel_tmp31_fu_1398_p2 = (working_key[3221] == 1'b1)? tmp75_fu_1393_p2 >> icmp_ln123_reg_4642 : tmp75_fu_1393_p2 & icmp_ln123_reg_4642;
  assign sel_tmp37_fu_1403_p2 = (working_key[3222] == 1'b1)? xor_ln118_fu_1377_p2 & icmp_ln123_2_reg_4668 : xor_ln118_fu_1377_p2 | icmp_ln123_2_reg_4668;
  assign sel_tmp50_fu_2293_p2 = (working_key[3223] == 1'b1)? tmp110_fu_2287_p2 ^ icmp_ln123_4_fu_2219_p2 : tmp110_fu_2287_p2 & icmp_ln123_4_fu_2219_p2;
  assign sel_tmp57_fu_2321_p2 = (working_key[3224] == 1'b1)? tmp111_fu_2315_p2 & icmp_ln123_3_fu_2203_p2 : tmp111_fu_2315_p2 ^ icmp_ln123_3_fu_2203_p2;
  assign sel_tmp63_fu_2343_p2 = (working_key[3225] == 1'b1)? xor_ln118_1_fu_2281_p2 >> icmp_ln123_6_fu_2337_p2 : xor_ln118_1_fu_2281_p2 & icmp_ln123_6_fu_2337_p2;
  assign Const_978 = (1'd0 ^ working_key[3226]);
  assign Const_979 = (24'd5854932 ^ working_key[3251:3228]);
  assign Const_980 = (24'd5396139 ^ working_key[3275:3252]);
  assign select_ln116_1_fu_1173_p3 = ((((working_key[3227] == 1'b1)? tmp_1_fu_1157_p3[0:0] != Const_978 : tmp_1_fu_1157_p3[0:0] === Const_978) ^ working_key[3276]) == 1'b1)? Const_980 : Const_979;
  assign Const_981 = (1'd1 ^ working_key[3277]);
  assign Const_982 = (32'd2863484950 ^ working_key[3310:3279]);
  assign Const_983 = (32'd1431654485 ^ working_key[3342:3311]);
  assign select_ln116_2_fu_2121_p3 = ((((working_key[3278] == 1'b1)? tmp_16_fu_2113_p3[0:0] === Const_981 : tmp_16_fu_2113_p3[0:0] < Const_981) ^ working_key[3343]) == 1'b1)? Const_983 : Const_982;
  assign Const_984 = (1'd1 ^ working_key[3344]);
  assign Const_985 = (24'd5984900 ^ working_key[3369:3346]);
  assign Const_986 = (24'd5942938 ^ working_key[3393:3370]);
  assign select_ln116_3_fu_2133_p3 = ((((working_key[3345] == 1'b1)? tmp_16_fu_2113_p3[0:0] > Const_984 : tmp_16_fu_2113_p3[0:0] === Const_984) ^ working_key[3394]) == 1'b1)? Const_986 : Const_985;
  assign Const_987 = (1'd1 ^ working_key[3395]);
  assign Const_988 = (16'd22870 ^ working_key[3412:3397]);
  assign Const_989 = (16'd19135 ^ working_key[3428:3413]);
  assign select_ln116_4_fu_2145_p3 = ((((working_key[3396] == 1'b1)? tmp_16_fu_2113_p3[0:0] != Const_987 : tmp_16_fu_2113_p3[0:0] === Const_987) ^ working_key[3429]) == 1'b1)? Const_989 : Const_988;
  assign Const_990 = (1'd1 ^ working_key[3430]);
  assign Const_991 = (8'd85 ^ working_key[3439:3432]);
  assign Const_992 = (8'd42 ^ working_key[3447:3440]);
  assign select_ln116_5_fu_2157_p3 = ((((working_key[3431] == 1'b1)? tmp_16_fu_2113_p3[0:0] === Const_990 : tmp_16_fu_2113_p3[0:0] < Const_990) ^ working_key[3448]) == 1'b1)? Const_991 : Const_992;
  assign Const_993 = (1'd1 ^ working_key[3449]);
  assign Const_994 = (32'd1449831082 ^ working_key[3482:3451]);
  assign Const_995 = (32'd1464685142 ^ working_key[3514:3483]);
  assign select_ln116_fu_1165_p3 = ((((working_key[3450] == 1'b1)? tmp_1_fu_1157_p3[0:0] != Const_993 : tmp_1_fu_1157_p3[0:0] === Const_993) ^ working_key[3515]) == 1'b1)? Const_995 : Const_994;
  assign Const_996 = (1'd1 ^ working_key[3516]);
  assign select_ln118_1_fu_2414_p3 = ((((working_key[3517] == 1'b1)? sel_tmp57_reg_5277[0:0] === Const_996 : sel_tmp57_reg_5277[0:0] == Const_996) ^ working_key[3518]) == 1'b1)? zext_ln123_9_fu_2393_p1 : add_ln123_3_fu_2381_p2;
  assign Const_997 = (1'd1 ^ working_key[3519]);
  assign select_ln118_2_fu_2421_p3 = ((((working_key[3520] == 1'b1)? or_ln118_reg_5282[0:0] === Const_997 : or_ln118_reg_5282[0:0] < Const_997) ^ working_key[3521]) == 1'b1)? select_ln118_fu_2407_p3 : select_ln118_1_fu_2414_p3;
  assign Const_998 = (1'd0 ^ working_key[3522]);
  assign Const_999 = (5'd18 ^ working_key[3528:3524]);
  assign select_ln118_fu_2407_p3 = ((((working_key[3523] == 1'b1)? icmp_ln118_1_reg_5252[0:0] == Const_998 : icmp_ln118_1_reg_5252[0:0] === Const_998) ^ working_key[3529]) == 1'b1)? Const_999 : add_ln123_2_fu_2371_p2;
  assign Const_1000 = (1'd0 ^ working_key[3530]);
  assign Const_1001 = (64'd12297785402006536114 ^ working_key[3595:3532]);
  assign Const_1002 = (64'd2696172293825363658 ^ working_key[3659:3596]);
  assign select_ln123_fu_1237_p3 = ((((working_key[3531] == 1'b1)? tmp_1_fu_1157_p3[0:0] == Const_1000 : tmp_1_fu_1157_p3[0:0] === Const_1000) ^ working_key[3660]) == 1'b1)? Const_1002 : Const_1001;
  assign Const_1003 = (1'd1 ^ working_key[3661]);
  assign select_ln213_fu_2648_p3 = ((((working_key[3662] == 1'b1)? icmp_ln213_fu_2637_p2[0:0] === Const_1003 : icmp_ln213_fu_2637_p2[0:0] > Const_1003) ^ working_key[3663]) == 1'b1)? sub_ln214_fu_2642_p2 : ap_phi_mux_p_0_i52_i_phi_fu_1041_p4;
  assign Const_1004 = (1'd0 ^ working_key[3664]);
  assign select_ln273_fu_3151_p3 = ((((working_key[3665] == 1'b1)? tmp_39_fu_3037_p3[0:0] != Const_1004 : tmp_39_fu_3037_p3[0:0] === Const_1004) ^ working_key[3666]) == 1'b1)? temp_23_fu_3137_p3 : sub_ln273_fu_3145_p2;
  assign Const_1005 = (1'd0 ^ working_key[3667]);
  assign select_ln304_1_fu_3654_p3 = ((((working_key[3668] == 1'b1)? or_ln304_fu_3648_p2[0:0] == Const_1005 : or_ln304_fu_3648_p2[0:0] === Const_1005) ^ working_key[3669]) == 1'b1)? select_ln304_fu_3640_p3 : add_ln304_fu_3634_p2;
  assign Const_1006 = (1'd0 ^ working_key[3670]);
  assign Const_1007 = (8'd64 ^ working_key[3679:3672]);
  assign Const_1008 = (8'd149 ^ working_key[3687:3680]);
  assign select_ln304_fu_3640_p3 = ((((working_key[3671] == 1'b1)? icmp_ln304_fu_3622_p2[0:0] < Const_1006 : icmp_ln304_fu_3622_p2[0:0] === Const_1006) ^ working_key[3688]) == 1'b1)? Const_1007 : Const_1008;
  assign Const_1009 = (1'd0 ^ working_key[3689]);
  assign select_ln305_1_fu_3719_p3 = ((((working_key[3690] == 1'b1)? or_ln305_fu_3713_p2[0:0] != Const_1009 : or_ln305_fu_3713_p2[0:0] === Const_1009) ^ working_key[3691]) == 1'b1)? add_ln305_fu_3699_p2 : select_ln305_fu_3705_p3;
  assign Const_1010 = (1'd1 ^ working_key[3692]);
  assign Const_1011 = (8'd149 ^ working_key[3701:3694]);
  assign Const_1012 = (8'd10 ^ working_key[3709:3702]);
  assign select_ln305_fu_3705_p3 = ((((working_key[3693] == 1'b1)? icmp_ln305_fu_3687_p2[0:0] === Const_1010 : icmp_ln305_fu_3687_p2[0:0] == Const_1010) ^ working_key[3710]) == 1'b1)? Const_1011 : Const_1012;
  assign Const_1013 = (1'd0 ^ working_key[3711]);
  assign select_ln306_1_fu_3890_p3 = ((((working_key[3712] == 1'b1)? or_ln306_fu_3884_p2[0:0] == Const_1013 : or_ln306_fu_3884_p2[0:0] === Const_1013) ^ working_key[3713]) == 1'b1)? add_ln306_fu_3870_p2 : select_ln306_fu_3876_p3;
  assign Const_1014 = (1'd1 ^ working_key[3714]);
  assign Const_1015 = (8'd181 ^ working_key[3723:3716]);
  assign Const_1016 = (8'd170 ^ working_key[3731:3724]);
  assign select_ln306_fu_3876_p3 = ((((working_key[3715] == 1'b1)? icmp_ln306_fu_3858_p2[0:0] === Const_1014 : icmp_ln306_fu_3858_p2[0:0] > Const_1014) ^ working_key[3732]) == 1'b1)? Const_1015 : Const_1016;
  assign Const_1017 = (1'd1 ^ working_key[3733]);
  assign select_ln307_1_fu_3955_p3 = ((((working_key[3734] == 1'b1)? or_ln307_fu_3949_p2[0:0] === Const_1017 : or_ln307_fu_3949_p2[0:0] != Const_1017) ^ working_key[3735]) == 1'b1)? add_ln307_fu_3935_p2 : select_ln307_fu_3941_p3;
  assign Const_1018 = (1'd1 ^ working_key[3736]);
  assign Const_1019 = (8'd202 ^ working_key[3745:3738]);
  assign Const_1020 = (8'd74 ^ working_key[3753:3746]);
  assign select_ln307_fu_3941_p3 = ((((working_key[3737] == 1'b1)? icmp_ln307_fu_3923_p2[0:0] < Const_1018 : icmp_ln307_fu_3923_p2[0:0] === Const_1018) ^ working_key[3754]) == 1'b1)? Const_1019 : Const_1020;
  assign Const_1021 = (1'd0 ^ working_key[3755]);
  assign select_ln309_1_fu_4080_p3 = ((((working_key[3756] == 1'b1)? or_ln309_fu_4074_p2[0:0] == Const_1021 : or_ln309_fu_4074_p2[0:0] === Const_1021) ^ working_key[3757]) == 1'b1)? add_ln309_fu_4060_p2 : select_ln309_fu_4066_p3;
  assign Const_1022 = (1'd1 ^ working_key[3758]);
  assign Const_1023 = (8'd169 ^ working_key[3767:3760]);
  assign Const_1024 = (8'd171 ^ working_key[3775:3768]);
  assign select_ln309_fu_4066_p3 = ((((working_key[3759] == 1'b1)? icmp_ln309_fu_4048_p2[0:0] === Const_1022 : icmp_ln309_fu_4048_p2[0:0] == Const_1022) ^ working_key[3776]) == 1'b1)? Const_1023 : Const_1024;
  assign Const_1025 = (1'd0 ^ working_key[3777]);
  assign select_ln310_1_fu_4145_p3 = ((((working_key[3778] == 1'b1)? or_ln310_fu_4139_p2[0:0] === Const_1025 : or_ln310_fu_4139_p2[0:0] > Const_1025) ^ working_key[3779]) == 1'b1)? select_ln310_fu_4131_p3 : add_ln310_fu_4125_p2;
  assign Const_1026 = (1'd0 ^ working_key[3780]);
  assign Const_1027 = (8'd70 ^ working_key[3789:3782]);
  assign Const_1028 = (8'd53 ^ working_key[3797:3790]);
  assign select_ln310_fu_4131_p3 = ((((working_key[3781] == 1'b1)? icmp_ln310_fu_4113_p2[0:0] == Const_1026 : icmp_ln310_fu_4113_p2[0:0] === Const_1026) ^ working_key[3798]) == 1'b1)? Const_1028 : Const_1027;
  assign Const_1029 = (1'd1 ^ working_key[3799]);
  assign select_ln311_1_fu_4210_p3 = ((((working_key[3800] == 1'b1)? or_ln311_fu_4204_p2[0:0] === Const_1029 : or_ln311_fu_4204_p2[0:0] != Const_1029) ^ working_key[3801]) == 1'b1)? add_ln311_fu_4190_p2 : select_ln311_fu_4196_p3;
  assign Const_1030 = (1'd0 ^ working_key[3802]);
  assign Const_1031 = (8'd80 ^ working_key[3811:3804]);
  assign Const_1032 = (8'd169 ^ working_key[3819:3812]);
  assign select_ln311_fu_4196_p3 = ((((working_key[3803] == 1'b1)? icmp_ln311_fu_4178_p2[0:0] === Const_1030 : icmp_ln311_fu_4178_p2[0:0] != Const_1030) ^ working_key[3820]) == 1'b1)? Const_1031 : Const_1032;
  assign Const_1033 = (1'd0 ^ working_key[3821]);
  assign select_ln312_1_fu_4275_p3 = ((((working_key[3822] == 1'b1)? or_ln312_fu_4269_p2[0:0] != Const_1033 : or_ln312_fu_4269_p2[0:0] === Const_1033) ^ working_key[3823]) == 1'b1)? add_ln312_fu_4255_p2 : select_ln312_fu_4261_p3;
  assign Const_1034 = (1'd1 ^ working_key[3824]);
  assign Const_1035 = (8'd173 ^ working_key[3833:3826]);
  assign Const_1036 = (8'd160 ^ working_key[3841:3834]);
  assign select_ln312_fu_4261_p3 = ((((working_key[3825] == 1'b1)? icmp_ln312_fu_4243_p2[0:0] === Const_1034 : icmp_ln312_fu_4243_p2[0:0] > Const_1034) ^ working_key[3842]) == 1'b1)? Const_1035 : Const_1036;
  assign Const_1037 = (1'd0 ^ working_key[3843]);
  assign Const_1038 = (7'd21 ^ working_key[3851:3845]);
  assign select_ln40_10_fu_3903_p3 = ((((working_key[3844] == 1'b1)? icmp_ln40_8_reg_5597[0:0] > Const_1037 : icmp_ln40_8_reg_5597[0:0] === Const_1037) ^ working_key[3852]) == 1'b1)? Const_1038 : tmp_8_reg_5602;
  assign Const_1039 = (1'd0 ^ working_key[3853]);
  assign Const_1040 = (7'd42 ^ working_key[3861:3855]);
  assign select_ln40_12_fu_4028_p3 = ((((working_key[3854] == 1'b1)? icmp_ln40_12_reg_5643[0:0] < Const_1039 : icmp_ln40_12_reg_5643[0:0] === Const_1039) ^ working_key[3862]) == 1'b1)? tmp_9_reg_5648 : Const_1040;
  assign Const_1041 = (1'd0 ^ working_key[3863]);
  assign Const_1042 = (7'd111 ^ working_key[3871:3865]);
  assign select_ln40_13_fu_4093_p3 = ((((working_key[3864] == 1'b1)? icmp_ln40_13_reg_5623[0:0] > Const_1041 : icmp_ln40_13_reg_5623[0:0] === Const_1041) ^ working_key[3872]) == 1'b1)? tmp_s_reg_5628 : Const_1042;
  assign Const_1043 = (1'd0 ^ working_key[3873]);
  assign Const_1044 = (7'd101 ^ working_key[3881:3875]);
  assign select_ln40_14_fu_4158_p3 = ((((working_key[3874] == 1'b1)? icmp_ln40_14_reg_5665[0:0] < Const_1043 : icmp_ln40_14_reg_5665[0:0] === Const_1043) ^ working_key[3882]) == 1'b1)? Const_1044 : tmp_10_reg_5670;
  assign Const_1045 = (1'd0 ^ working_key[3883]);
  assign Const_1046 = (7'd117 ^ working_key[3891:3885]);
  assign select_ln40_15_fu_4223_p3 = ((((working_key[3884] == 1'b1)? icmp_ln40_15_reg_5675[0:0] == Const_1045 : icmp_ln40_15_reg_5675[0:0] === Const_1045) ^ working_key[3892]) == 1'b1)? Const_1046 : tmp_11_reg_5680;
  assign Const_1047 = (1'd0 ^ working_key[3893]);
  assign select_ln40_1_fu_2774_p3 = ((((working_key[3894] == 1'b1)? or_ln40_fu_2768_p2[0:0] < Const_1047 : or_ln40_fu_2768_p2[0:0] === Const_1047) ^ working_key[3895]) == 1'b1)? add_ln40_1_fu_2754_p2 : select_ln40_fu_2760_p3;
  assign Const_1048 = (1'd0 ^ working_key[3896]);
  assign Const_1049 = (16'd5546 ^ working_key[3913:3898]);
  assign Const_1050 = (16'd44203 ^ working_key[3929:3914]);
  assign select_ln40_2_fu_2922_p3 = ((((working_key[3897] == 1'b1)? icmp_ln40_2_fu_2895_p2[0:0] === Const_1048 : icmp_ln40_2_fu_2895_p2[0:0] == Const_1048) ^ working_key[3930]) == 1'b1)? Const_1050 : Const_1049;
  assign Const_1051 = (1'd0 ^ working_key[3931]);
  assign select_ln40_3_fu_2936_p3 = ((((working_key[3932] == 1'b1)? or_ln40_1_fu_2930_p2[0:0] === Const_1051 : or_ln40_1_fu_2930_p2[0:0] > Const_1051) ^ working_key[3933]) == 1'b1)? add_ln40_6_fu_2917_p2 : select_ln40_2_fu_2922_p3;
  assign Const_1052 = (1'd0 ^ working_key[3934]);
  assign Const_1053 = (16'd10901 ^ working_key[3951:3936]);
  assign Const_1054 = (16'd64853 ^ working_key[3967:3952]);
  assign select_ln40_4_fu_2980_p3 = ((((working_key[3935] == 1'b1)? icmp_ln40_4_fu_2954_p2[0:0] == Const_1052 : icmp_ln40_4_fu_2954_p2[0:0] === Const_1052) ^ working_key[3968]) == 1'b1)? Const_1053 : Const_1054;
  assign Const_1055 = (1'd0 ^ working_key[3969]);
  assign select_ln40_5_fu_2994_p3 = ((((working_key[3970] == 1'b1)? or_ln40_2_fu_2988_p2[0:0] != Const_1055 : or_ln40_2_fu_2988_p2[0:0] === Const_1055) ^ working_key[3971]) == 1'b1)? add_ln40_10_fu_2976_p2 : select_ln40_4_fu_2980_p3;
  assign Const_1056 = (1'd1 ^ working_key[3972]);
  assign Const_1057 = (7'd21 ^ working_key[3980:3974]);
  assign select_ln40_6_fu_3602_p3 = ((((working_key[3973] == 1'b1)? icmp_ln40_6_reg_5557[0:0] === Const_1056 : icmp_ln40_6_reg_5557[0:0] != Const_1056) ^ working_key[3981]) == 1'b1)? tmp_5_reg_5562 : Const_1057;
  assign Const_1058 = (1'd1 ^ working_key[3982]);
  assign Const_1059 = (7'd117 ^ working_key[3990:3984]);
  assign select_ln40_7_fu_3667_p3 = ((((working_key[3983] == 1'b1)? icmp_ln40_7_reg_5567[0:0] === Const_1058 : icmp_ln40_7_reg_5567[0:0] == Const_1058) ^ working_key[3991]) == 1'b1)? tmp_6_reg_5572 : Const_1059;
  assign Const_1060 = (1'd1 ^ working_key[3992]);
  assign Const_1061 = (7'd106 ^ working_key[4000:3994]);
  assign select_ln40_9_fu_3838_p3 = ((((working_key[3993] == 1'b1)? icmp_ln40_10_reg_5587[0:0] != Const_1060 : icmp_ln40_10_reg_5587[0:0] === Const_1060) ^ working_key[4001]) == 1'b1)? tmp_7_reg_5592 : Const_1061;
  assign Const_1062 = (1'd1 ^ working_key[4002]);
  assign Const_1063 = (16'd60050 ^ working_key[4019:4004]);
  assign Const_1064 = (16'd5445 ^ working_key[4035:4020]);
  assign select_ln40_fu_2760_p3 = ((((working_key[4003] == 1'b1)? icmp_ln40_fu_2732_p2[0:0] === Const_1062 : icmp_ln40_fu_2732_p2[0:0] != Const_1062) ^ working_key[4036]) == 1'b1)? Const_1064 : Const_1063;
  assign Const_1065 = (1'd1 ^ working_key[4037]);
  assign select_ln61_fu_1334_p3 = ((((working_key[4038] == 1'b1)? icmp_ln61_fu_1328_p2[0:0] === Const_1065 : icmp_ln61_fu_1328_p2[0:0] > Const_1065) ^ working_key[4039]) == 1'b1)? smax_fu_1320_p3 : smax_0_i_reg_839;
  assign Const_1066 = (1'd1 ^ working_key[4040]);
  assign Const_1067 = (6'd20 ^ working_key[4047:4042]);
  assign Const_1068 = (6'd9 ^ working_key[4053:4048]);
  assign select_ln67_fu_1458_p3 = ((((working_key[4041] == 1'b1)? icmp_ln67_fu_1342_p2[0:0] === Const_1066 : icmp_ln67_fu_1342_p2[0:0] != Const_1066) ^ working_key[4054]) == 1'b1)? Const_1068 : Const_1067;
  assign Const_1069 = (1'd1 ^ working_key[4055]);
  assign Const_1070 = (15'd13632 ^ working_key[4071:4057]);
  assign select_ln72_1_fu_2543_p3 = ((((working_key[4056] == 1'b1)? grp_fu_1093_p2[0:0] === Const_1069 : grp_fu_1093_p2[0:0] > Const_1069) ^ working_key[4072]) == 1'b1)? Const_1070 : sub_ln72_1_fu_2537_p2;
  assign Const_1071 = (1'd0 ^ working_key[4073]);
  assign Const_1072 = (16'd10922 ^ working_key[4090:4075]);
  assign select_ln72_2_fu_3057_p3 = ((((working_key[4074] == 1'b1)? icmp_ln72_4_fu_3045_p2[0:0] != Const_1071 : icmp_ln72_4_fu_3045_p2[0:0] === Const_1071) ^ working_key[4091]) == 1'b1)? Const_1072 : sub_ln72_2_fu_3051_p2;
  assign Const_1073 = (1'd1 ^ working_key[4092]);
  assign Const_1074 = (16'd54613 ^ working_key[4109:4094]);
  assign select_ln72_fu_1312_p3 = ((((working_key[4093] == 1'b1)? icmp_ln72_1_fu_1300_p2[0:0] == Const_1073 : icmp_ln72_1_fu_1300_p2[0:0] === Const_1073) ^ working_key[4110]) == 1'b1)? Const_1074 : sub_ln72_fu_1306_p2;
  assign sext_ln100_1_fu_1596_p1 = sl_3_reg_4760;
  assign sext_ln100_fu_1593_p1 = sl_3_reg_4760;
  assign sext_ln105_1_fu_1599_p1 = sl_4_reg_4788;
  assign sext_ln109_fu_1751_p1 = mul_ln109_reg_4957;
  assign sext_ln111_1_fu_1605_p1 = sl_5_reg_4794;
  assign sext_ln111_2_fu_1754_p1 = mul_ln111_reg_4962;
  assign sext_ln111_fu_1602_p1 = sl_5_reg_4794;
  assign sext_ln116_fu_1641_p1 = mul_ln116_reg_4906;
  assign sext_ln118_1_fu_1612_p0 = s_q1;
  assign sext_ln118_1_fu_1612_p1 = sext_ln118_1_fu_1612_p0;
  assign sext_ln123_2_fu_2403_p1 = add_ln123_5_fu_2397_p2;
  assign sext_ln123_fu_1368_p1 = add_ln123_1_fu_1362_p2;
  assign sext_ln126_1_fu_1662_p0 = reg_1099;
  assign sext_ln126_1_fu_1662_p1 = sext_ln126_1_fu_1662_p0;
  assign sext_ln126_3_fu_1763_p1 = add_ln126_2_reg_4973;
  assign sext_ln126_4_fu_1666_p1 = grp_fu_4390_p3;
  assign sext_ln126_5_fu_1669_p1 = grp_fu_4397_p3;
  assign sext_ln126_6_fu_1772_p1 = add_ln126_7_reg_4978;
  assign sext_ln127_1_fu_1684_p1 = mul_ln127_reg_4947;
  assign sext_ln127_6_fu_1696_p1 = grp_fu_4456_p4;
  assign sext_ln128_1_fu_1705_p1 = grp_fu_4403_p3;
  assign sext_ln128_2_fu_1714_p1 = grp_fu_4430_p3;
  assign sext_ln128_3_fu_1717_p1 = grp_fu_4465_p3;
  assign sext_ln128_4_fu_1726_p1 = add_ln128_5_fu_1720_p2;
  assign sext_ln129_1_fu_1782_p1 = add_ln129_1_reg_4993;
  assign sext_ln129_2_fu_1791_p1 = add_ln129_4_reg_4998;
  assign sext_ln130_1_fu_1806_p1 = add_ln130_3_reg_5003;
  assign sext_ln131_1_fu_1742_p1 = grp_fu_4489_p3;
  assign sext_ln132_1_fu_1815_p1 = add_ln132_1_reg_5013;
  assign sext_ln133_fu_1824_p1 = mul_ln133_reg_5018;
  assign sext_ln138_fu_2561_p1 = temp_24_reg_997;
  assign sext_ln139_1_fu_2569_p0 = P_q0;
  assign sext_ln139_1_fu_2569_p1 = sext_ln139_1_fu_2569_p0;
  assign sext_ln139_fu_2565_p0 = P_q0;
  assign sext_ln139_fu_2565_p1 = sext_ln139_fu_2565_p0;
  assign sext_ln140_1_fu_1968_p1 = mul_ln140_reg_5121;
  assign sext_ln140_fu_1882_p1 = reg_1099;
  assign sext_ln141_1_fu_1916_p1 = mul_ln141_reg_5101;
  assign sext_ln142_1_fu_1925_p1 = mul_ln142_reg_5106;
  assign sext_ln143_1_fu_1978_p1 = mul_ln143_reg_5136;
  assign sext_ln144_1_fu_1987_p1 = mul_ln144_reg_5141;
  assign sext_ln145_1_fu_2004_p1 = mul_ln145_reg_5171;
  assign sext_ln146_1_fu_2013_p1 = mul_ln146_reg_5176;
  assign sext_ln147_1_fu_2030_p1 = mul_ln147_reg_5201;
  assign sext_ln148_1_fu_2039_p1 = mul_ln148_reg_5206;
  assign sext_ln151_fu_2048_p1 = k_3_i_reg_906;
  assign sext_ln187_fu_2439_p1 = temp_2_fu_2432_p3;
  assign sext_ln304_1_fu_3662_p1 = select_ln304_1_fu_3654_p3;
  assign sext_ln304_fu_3608_p1 = select_ln40_6_fu_3602_p3;
  assign sext_ln305_1_fu_3727_p1 = select_ln305_1_fu_3719_p3;
  assign sext_ln305_fu_3673_p1 = select_ln40_7_fu_3667_p3;
  assign sext_ln306_1_fu_3898_p1 = select_ln306_1_fu_3890_p3;
  assign sext_ln306_fu_3844_p1 = select_ln40_9_fu_3838_p3;
  assign sext_ln307_1_fu_3963_p1 = select_ln307_1_fu_3955_p3;
  assign sext_ln307_fu_3909_p1 = select_ln40_10_fu_3903_p3;
  assign sext_ln309_1_fu_4088_p1 = select_ln309_1_fu_4080_p3;
  assign sext_ln309_fu_4034_p1 = select_ln40_12_fu_4028_p3;
  assign sext_ln310_1_fu_4153_p1 = select_ln310_1_fu_4145_p3;
  assign sext_ln310_fu_4099_p1 = select_ln40_13_fu_4093_p3;
  assign sext_ln311_1_fu_4218_p1 = select_ln311_1_fu_4210_p3;
  assign sext_ln311_fu_4164_p1 = select_ln40_14_fu_4158_p3;
  assign sext_ln312_1_fu_4283_p1 = select_ln312_1_fu_4275_p3;
  assign sext_ln312_fu_4229_p1 = select_ln40_15_fu_4223_p3;
  assign sext_ln39_10_fu_3732_p1 = temp_13_reg_5617;
  assign sext_ln39_11_fu_3770_p1 = temp_14_fu_3762_p3;
  assign sext_ln39_12_fu_3570_p1 = temp_15_fu_3560_p4;
  assign sext_ln39_13_fu_3968_p1 = temp_16_reg_5653;
  assign sext_ln39_14_fu_3998_p1 = temp_17_reg_5659;
  assign sext_ln39_2_fu_2882_p1 = reg_1122;
  assign sext_ln39_3_fu_2886_p1 = temp_6_reg_5512;
  assign sext_ln39_4_fu_2945_p1 = temp_7_reg_5518;
  assign sext_ln39_5_fu_3199_p1 = temp_8_fu_3189_p4;
  assign sext_ln39_6_fu_3281_p1 = temp_9_fu_3271_p4;
  assign sext_ln39_7_fu_3363_p1 = temp_10_fu_3353_p4;
  assign sext_ln39_8_fu_3403_p1 = temp_11_fu_3395_p3;
  assign sext_ln39_9_fu_3485_p1 = temp_12_fu_3475_p4;
  assign sext_ln39_fu_2723_p1 = temp_5_fu_2715_p3;
  assign sext_ln50_10_fu_3550_p1 = shl_ln50_9_fu_3542_p3;
  assign sext_ln50_1_fu_3179_p1 = shl_ln50_1_fu_3171_p3;
  assign sext_ln50_2_fu_3249_p1 = shl_ln50_2_fu_3241_p3;
  assign sext_ln50_3_fu_3261_p1 = shl_ln50_3_fu_3253_p3;
  assign sext_ln50_4_fu_3331_p1 = shl_ln50_4_fu_3323_p3;
  assign sext_ln50_5_fu_3343_p1 = shl_ln50_5_fu_3335_p3;
  assign sext_ln50_6_fu_3453_p1 = shl_ln50_6_fu_3445_p3;
  assign sext_ln50_7_fu_3465_p1 = shl_ln50_7_fu_3457_p3;
  assign sext_ln50_9_fu_3538_p1 = shl_ln50_8_fu_3530_p3;
  assign sext_ln50_fu_3167_p1 = shl_ln1_fu_3159_p3;
  assign sext_ln62_2_fu_2703_p1 = select_ln213_reg_5434;
  assign sext_ln62_3_fu_2879_p1 = K_load_reg_5506;
  assign sext_ln67_fu_1479_p1 = n_fu_1471_p3;
  assign sext_ln88_fu_1554_p1 = k_2_i_reg_873;
  assign sext_ln91_fu_1577_p1 = reg_1099;
  assign sext_ln93_1_fu_1584_p1 = sl_1_reg_4732;
  assign sext_ln94_fu_1623_p1 = mul_ln94_reg_4831;
  assign sext_ln96_1_fu_1590_p1 = sl_2_reg_4754;
  assign Const_1075 = (64'd12270854832493259156 ^ working_key[4174:4111]);
  assign shl_ln152_fu_2071_p2 = (working_key[4175] == 1'b1)? L_ACF_q0 << Const_1075 : L_ACF_q0 >> Const_1075;
  assign shl_ln187_fu_2464_p2 = (working_key[4176] == 1'b1)? trunc_ln187_fu_2460_p1 >> sext_ln187_reg_5292 : trunc_ln187_fu_2460_p1 << sext_ln187_reg_5292;
  assign shl_ln1_fu_3159_p3 = { { LARc_q0 }, { 14'd0 } };
  assign Const_1076 = (16'd44024 ^ working_key[4192:4177]);
  assign shl_ln270_fu_3105_p2 = (working_key[4193] == 1'b1)? temp_fu_3065_p3 >> Const_1076 : temp_fu_3065_p3 << Const_1076;
  assign shl_ln50_1_fu_3171_p3 = { { LARc_q0 }, { 12'd0 } };
  assign shl_ln50_2_fu_3241_p3 = { { LARc_q1 }, { 14'd0 } };
  assign shl_ln50_3_fu_3253_p3 = { { LARc_q1 }, { 12'd0 } };
  assign shl_ln50_4_fu_3323_p3 = { { LARc_q1 }, { 14'd0 } };
  assign shl_ln50_5_fu_3335_p3 = { { LARc_q1 }, { 12'd0 } };
  assign shl_ln50_6_fu_3445_p3 = { { LARc_q0 }, { 14'd0 } };
  assign shl_ln50_7_fu_3457_p3 = { { LARc_q0 }, { 12'd0 } };
  assign shl_ln50_8_fu_3530_p3 = { { LARc_q0 }, { 14'd0 } };
  assign shl_ln50_9_fu_3542_p3 = { { LARc_q0 }, { 10'd0 } };
  assign Const_1077 = (1'd1 ^ working_key[4194]);
  assign smax_fu_1320_p3 = ((((working_key[4195] == 1'b1)? tmp_13_fu_1292_p3[0:0] === Const_1077 : tmp_13_fu_1292_p3[0:0] == Const_1077) ^ working_key[4196]) == 1'b1)? select_ln72_fu_1312_p3 : s_q0;
  assign sp_0_rec_i_cast_fu_1833_p1 = sp_0_rec_i_reg_894;
  assign Const_1078 = (16'd21845 ^ working_key[4212:4197]);
  assign sub_ln214_fu_2642_p2 = (working_key[4213] == 1'b1)? Const_1078 - ap_phi_mux_p_0_i52_i_phi_fu_1041_p4 : Const_1078 << ap_phi_mux_p_0_i52_i_phi_fu_1041_p4;
  assign Const_1079 = (32'd850045608 ^ working_key[4245:4214]);
  assign sub_ln223_fu_2782_p2 = (working_key[4246] == 1'b1)? Const_1079 - i_3_reg_973 : Const_1079 * i_3_reg_973;
  assign Const_1080 = (16'd9578 ^ working_key[4262:4247]);
  assign sub_ln273_fu_3145_p2 = (working_key[4263] == 1'b1)? Const_1080 - temp_23_fu_3137_p3 : Const_1080 * temp_23_fu_3137_p3;
  assign sub_ln50_fu_3554_p2 = (working_key[4264] == 1'b1)? sext_ln50_9_fu_3538_p1 * sext_ln50_10_fu_3550_p1 : sext_ln50_9_fu_3538_p1 - sext_ln50_10_fu_3550_p1;
  assign Const_1081 = (6'd49 ^ working_key[4270:4265]);
  assign sub_ln70_fu_1452_p2 = (working_key[4271] == 1'b1)? Const_1081 << newSel114_fu_1444_p3 : Const_1081 - newSel114_fu_1444_p3;
  assign Const_1082 = (15'd27322 ^ working_key[4286:4272]);
  assign sub_ln72_1_fu_2537_p2 = (working_key[4287] == 1'b1)? Const_1082 + trunc_ln72_fu_2533_p1 : Const_1082 - trunc_ln72_fu_2533_p1;
  assign Const_1083 = (16'd54565 ^ working_key[4303:4288]);
  assign sub_ln72_2_fu_3051_p2 = (working_key[4304] == 1'b1)? Const_1083 + LARc_q0 : Const_1083 - LARc_q0;
  assign Const_1084 = (16'd44026 ^ working_key[4320:4305]);
  assign sub_ln72_fu_1306_p2 = (working_key[4321] == 1'b1)? Const_1084 * s_q0 : Const_1084 - s_q0;
  assign sum17_cast_fu_1843_p1 = sum17_fu_1837_p2;
  assign Const_1085 = (8'd173 ^ working_key[4329:4322]);
  assign sum17_fu_1837_p2 = (working_key[4330] == 1'b1)? sp_0_rec_i_reg_894 >> Const_1085 : sp_0_rec_i_reg_894 + Const_1085;
  assign sum42_cast_fu_2672_p1 = sum42_fu_2667_p2;
  assign sum42_fu_2667_p2 = (working_key[4331] == 1'b1)? empty_65_fu_2663_p1 + zext_ln206_1_reg_5411 : empty_65_fu_2663_p1 << zext_ln206_1_reg_5411;
  assign Const_1086 = (17'd97194 ^ working_key[4348:4332]);
  assign sum_10_fu_3574_p2 = (working_key[4349] == 1'b1)? sext_ln39_12_fu_3570_p1 + Const_1086 : sext_ln39_12_fu_3570_p1 * Const_1086;
  assign Const_1087 = (17'd87041 ^ working_key[4366:4350]);
  assign sum_11_fu_3971_p2 = (working_key[4367] == 1'b1)? sext_ln39_13_fu_3968_p1 + Const_1087 : sext_ln39_13_fu_3968_p1 << Const_1087;
  assign Const_1088 = (17'd85604 ^ working_key[4384:4368]);
  assign sum_12_fu_4001_p2 = (working_key[4385] == 1'b1)? sext_ln39_14_fu_3998_p1 + Const_1088 : sext_ln39_14_fu_3998_p1 >> Const_1088;
  assign sum_1_fu_2889_p2 = (working_key[4386] == 1'b1)? sext_ln39_2_fu_2882_p1 >> sext_ln39_3_fu_2886_p1 : sext_ln39_2_fu_2882_p1 + sext_ln39_3_fu_2886_p1;
  assign sum_2_fu_2948_p2 = (working_key[4387] == 1'b1)? sext_ln62_3_fu_2879_p1 << sext_ln39_4_fu_2945_p1 : sext_ln62_3_fu_2879_p1 + sext_ln39_4_fu_2945_p1;
  assign Const_1089 = (17'd108457 ^ working_key[4404:4388]);
  assign sum_3_fu_3203_p2 = (working_key[4405] == 1'b1)? sext_ln39_5_fu_3199_p1 + Const_1089 : sext_ln39_5_fu_3199_p1 * Const_1089;
  assign Const_1090 = (17'd38058 ^ working_key[4422:4406]);
  assign sum_4_fu_3285_p2 = (working_key[4423] == 1'b1)? sext_ln39_6_fu_3281_p1 >> Const_1090 : sext_ln39_6_fu_3281_p1 + Const_1090;
  assign Const_1091 = (17'd130261 ^ working_key[4440:4424]);
  assign sum_5_fu_3367_p2 = (working_key[4441] == 1'b1)? sext_ln39_7_fu_3363_p1 + Const_1091 : sext_ln39_7_fu_3363_p1 >> Const_1091;
  assign Const_1092 = (17'd43861 ^ working_key[4458:4442]);
  assign sum_6_fu_3407_p2 = (working_key[4459] == 1'b1)? sext_ln39_8_fu_3403_p1 + Const_1092 : sext_ln39_8_fu_3403_p1 << Const_1092;
  assign Const_1093 = (17'd95402 ^ working_key[4476:4460]);
  assign sum_7_fu_3489_p2 = (working_key[4477] == 1'b1)? sext_ln39_9_fu_3485_p1 + Const_1093 : sext_ln39_9_fu_3485_p1 >> Const_1093;
  assign Const_1094 = (17'd43764 ^ working_key[4494:4478]);
  assign sum_8_fu_3735_p2 = (working_key[4495] == 1'b1)? sext_ln39_10_fu_3732_p1 + Const_1094 : sext_ln39_10_fu_3732_p1 * Const_1094;
  assign Const_1095 = (17'd46156 ^ working_key[4512:4496]);
  assign sum_9_fu_3774_p2 = (working_key[4513] == 1'b1)? sext_ln39_11_fu_3770_p1 + Const_1095 : sext_ln39_11_fu_3770_p1 * Const_1095;
  assign sum_fu_2727_p2 = (working_key[4514] == 1'b1)? sext_ln139_1_reg_5402 * sext_ln39_fu_2723_p1 : sext_ln139_1_reg_5402 + sext_ln39_fu_2723_p1;
  assign temp_10_fu_3353_p4 = { { add_ln50_2_fu_3347_p2[30:15] } };
  assign Const_1096 = (1'd1 ^ working_key[4515]);
  assign Const_1097 = (16'd44203 ^ working_key[4532:4517]);
  assign temp_11_fu_3395_p3 = ((((working_key[4516] == 1'b1)? icmp_ln40_9_fu_3383_p2[0:0] === Const_1096 : icmp_ln40_9_fu_3383_p2[0:0] == Const_1096) ^ working_key[4533]) == 1'b1)? add_ln40_3_fu_3389_p2 : Const_1097;
  assign temp_12_fu_3475_p4 = { { add_ln50_3_fu_3469_p2[30:15] } };
  assign Const_1098 = (1'd1 ^ working_key[4534]);
  assign Const_1099 = (16'd23189 ^ working_key[4551:4536]);
  assign temp_14_fu_3762_p3 = ((((working_key[4535] == 1'b1)? icmp_ln40_11_fu_3751_p2[0:0] === Const_1098 : icmp_ln40_11_fu_3751_p2[0:0] != Const_1098) ^ working_key[4552]) == 1'b1)? add_ln40_7_fu_3757_p2 : Const_1099;
  assign temp_15_fu_3560_p4 = { { sub_ln50_fu_3554_p2[30:15] } };
  assign temp_19_fu_3089_p1 = trunc_ln5_fu_3079_p4;
  assign Const_1100 = (16'd11943 ^ working_key[4568:4553]);
  assign temp_20_fu_3099_p2 = (working_key[4569] == 1'b1)? Const_1100 + temp_fu_3065_p3 : Const_1100 - temp_fu_3065_p3;
  assign Const_1101 = (16'd49749 ^ working_key[4585:4570]);
  assign temp_21_fu_3111_p2 = (working_key[4586] == 1'b1)? Const_1101 * shl_ln270_fu_3105_p2 : Const_1101 + shl_ln270_fu_3105_p2;
  assign Const_1102 = (1'd0 ^ working_key[4587]);
  assign temp_22_fu_3117_p3 = ((((working_key[4588] == 1'b1)? icmp_ln259_fu_3073_p2[0:0] != Const_1102 : icmp_ln259_fu_3073_p2[0:0] === Const_1102) ^ working_key[4589]) == 1'b1)? temp_21_fu_3111_p2 : temp_19_fu_3089_p1;
  assign Const_1103 = (1'd1 ^ working_key[4590]);
  assign temp_23_fu_3137_p3 = ((((working_key[4591] == 1'b1)? and_ln263_fu_3131_p2[0:0] === Const_1103 : and_ln263_fu_3131_p2[0:0] < Const_1103) ^ working_key[4592]) == 1'b1)? temp_20_fu_3099_p2 : temp_22_fu_3117_p3;
  assign Const_1104 = (1'd0 ^ working_key[4593]);
  assign temp_2_fu_2432_p3 = ((((working_key[4594] == 1'b1)? or_ln118_2_reg_5287[0:0] == Const_1104 : or_ln118_2_reg_5287[0:0] === Const_1104) ^ working_key[4595]) == 1'b1)? sext_ln123_2_fu_2403_p1 : zext_ln118_fu_2428_p1;
  assign Const_1105 = (1'd1 ^ working_key[4596]);
  assign Const_1106 = (16'd54623 ^ working_key[4613:4598]);
  assign temp_5_fu_2715_p3 = ((((working_key[4597] == 1'b1)? and_ln58_fu_2694_p2[0:0] === Const_1105 : and_ln58_fu_2694_p2[0:0] < Const_1105) ^ working_key[4614]) == 1'b1)? Const_1106 : trunc_ln64_1_fu_2706_p4;
  assign Const_1107 = (1'd0 ^ working_key[4615]);
  assign Const_1108 = (16'd35242 ^ working_key[4632:4617]);
  assign temp_6_fu_2845_p3 = ((((working_key[4616] == 1'b1)? and_ln58_1_fu_2827_p2[0:0] > Const_1107 : and_ln58_1_fu_2827_p2[0:0] === Const_1107) ^ working_key[4633]) == 1'b1)? Const_1108 : trunc_ln64_2_fu_2836_p4;
  assign Const_1109 = (1'd0 ^ working_key[4634]);
  assign Const_1110 = (16'd54996 ^ working_key[4651:4636]);
  assign temp_7_fu_2871_p3 = ((((working_key[4635] == 1'b1)? and_ln58_2_fu_2857_p2[0:0] != Const_1109 : and_ln58_2_fu_2857_p2[0:0] === Const_1109) ^ working_key[4652]) == 1'b1)? Const_1110 : trunc_ln64_3_fu_2862_p4;
  assign temp_8_fu_3189_p4 = { { add_ln50_fu_3183_p2[30:15] } };
  assign temp_9_fu_3271_p4 = { { add_ln50_1_fu_3265_p2[30:15] } };
  assign Const_1111 = (1'd0 ^ working_key[4653]);
  assign temp_fu_3065_p3 = ((((working_key[4654] == 1'b1)? tmp_39_fu_3037_p3[0:0] === Const_1111 : tmp_39_fu_3037_p3[0:0] < Const_1111) ^ working_key[4655]) == 1'b1)? select_ln72_2_fu_3057_p3 : LARc_q0;
  assign tmp110_fu_2287_p2 = (working_key[4656] == 1'b1)? xor_ln123_1_fu_2275_p2 << xor_ln118_1_fu_2281_p2 : xor_ln123_1_fu_2275_p2 & xor_ln118_1_fu_2281_p2;
  assign tmp111_fu_2315_p2 = (working_key[4657] == 1'b1)? xor_ln118_1_fu_2281_p2 & icmp_ln123_5_fu_2309_p2 : xor_ln118_1_fu_2281_p2 | icmp_ln123_5_fu_2309_p2;
  assign tmp75_fu_1393_p2 = (working_key[4658] == 1'b1)? xor_ln118_fu_1377_p2 << tmp_1_reg_4637 : xor_ln118_fu_1377_p2 & tmp_1_reg_4637;
  assign tmp_13_fu_1292_p3 = s_q0[32'd15];
  assign tmp_14_fu_1558_p3 = k_2_i_reg_873[32'd4];
  assign tmp_15_fu_2052_p3 = k_3_i_reg_906[32'd4];
  assign tmp_16_fu_2113_p3 = L_ACF_q0[32'd63];
  assign tmp_17_fu_2193_p4 = { { xor_ln95_2_fu_2181_p2[31:16] } };
  assign tmp_18_fu_2209_p4 = { { xor_ln95_2_fu_2181_p2[31:24] } };
  assign tmp_19_fu_2299_p4 = { { xor_ln95_1_fu_2175_p2[15:8] } };
  assign tmp_1_fu_1157_p3 = smax_0_i_reg_839[32'd15];
  assign tmp_20_fu_2327_p4 = { { xor_ln95_2_fu_2181_p2[31:8] } };
  assign tmp_21_fu_2519_p1 = P_q0;
  assign tmp_21_fu_2519_p3 = tmp_21_fu_2519_p1[32'd15];
  assign tmp_22_fu_2738_p4 = { { sum_fu_2727_p2[16:15] } };
  assign tmp_23_fu_2901_p4 = { { sum_1_fu_2889_p2[16:15] } };
  assign tmp_24_fu_2960_p4 = { { sum_2_fu_2948_p2[16:15] } };
  assign tmp_25_fu_3209_p4 = { { sum_3_fu_3203_p2[16:15] } };
  assign tmp_26_fu_3612_p4 = { { select_ln40_6_fu_3602_p3[6:5] } };
  assign tmp_27_fu_3291_p4 = { { sum_4_fu_3285_p2[16:15] } };
  assign tmp_28_fu_3677_p4 = { { select_ln40_7_fu_3667_p3[6:5] } };
  assign tmp_29_fu_3373_p4 = { { sum_5_fu_3367_p2[16:15] } };
  assign tmp_2_fu_1205_p4 = { { xor_ln116_fu_1193_p2[31:16] } };
  assign tmp_30_fu_3413_p4 = { { sum_6_fu_3407_p2[16:15] } };
  assign tmp_31_fu_3848_p4 = { { select_ln40_9_fu_3838_p3[6:4] } };
  assign tmp_32_fu_3913_p4 = { { select_ln40_10_fu_3903_p3[6:4] } };
  assign tmp_33_fu_3741_p4 = { { sum_8_fu_3735_p2[16:15] } };
  assign tmp_34_fu_3780_p4 = { { sum_9_fu_3774_p2[16:15] } };
  assign tmp_35_fu_4038_p4 = { { select_ln40_12_fu_4028_p3[6:3] } };
  assign tmp_36_fu_4103_p4 = { { select_ln40_13_fu_4093_p3[6:3] } };
  assign tmp_37_fu_4168_p4 = { { select_ln40_14_fu_4158_p3[6:2] } };
  assign tmp_38_fu_4233_p4 = { { select_ln40_15_fu_4223_p3[6:2] } };
  assign tmp_39_fu_3037_p3 = LARc_q0[32'd15];
  assign tmp_3_fu_1221_p4 = { { xor_ln116_fu_1193_p2[31:24] } };
  assign tmp_4_fu_1276_p4 = { { xor_ln116_fu_1193_p2[31:8] } };
  assign tmp_fu_1382_p2 = (working_key[4659] == 1'b1)? xor_ln123_fu_1372_p2 & xor_ln118_fu_1377_p2 : xor_ln123_fu_1372_p2 | xor_ln118_fu_1377_p2;
  assign trunc_ln116_1_fu_1185_p3 = { { trunc_ln116_fu_1181_p1 }, { 16'd0 } };
  assign trunc_ln116_2_fu_2129_p1 = L_ACF_q0[31:0];
  assign trunc_ln116_3_fu_2141_p1 = L_ACF_q0[23:0];
  assign trunc_ln116_4_fu_2153_p1 = L_ACF_q0[15:0];
  assign trunc_ln116_5_fu_2165_p1 = L_ACF_q0[7:0];
  assign trunc_ln116_fu_1181_p1 = smax_0_i_reg_839[7:0];
  assign trunc_ln123_1_fu_1246_p4 = { { xor_ln116_1_fu_1199_p2[23:16] } };
  assign trunc_ln123_2_fu_1261_p4 = { { xor_ln116_fu_1193_p2[31:24] } };
  assign trunc_ln123_3_fu_2230_p4 = { { xor_ln95_1_fu_2175_p2[15:8] } };
  assign trunc_ln123_4_fu_2245_p4 = { { xor_ln95_3_fu_2187_p2[23:16] } };
  assign trunc_ln123_5_fu_2260_p4 = { { xor_ln95_2_fu_2181_p2[31:24] } };
  assign trunc_ln155_fu_2625_p1 = div_0_i_i_reg_1015[14:0];
  assign trunc_ln187_fu_2460_p1 = L_ACF_q1[31:0];
  assign trunc_ln5_fu_3079_p4 = { { temp_fu_3065_p3[15:1] } };
  assign trunc_ln64_1_fu_2706_p4 = { { grp_fu_4555_p3[30:15] } };
  assign trunc_ln64_2_fu_2836_p4 = { { grp_fu_4564_p3[30:15] } };
  assign trunc_ln64_3_fu_2862_p4 = { { grp_fu_4572_p3[30:15] } };
  assign trunc_ln72_fu_2533_p0 = P_q0;
  assign trunc_ln72_fu_2533_p1 = trunc_ln72_fu_2533_p0[14:0];
  assign trunc_ln76_fu_1501_p1 = n_fu_1471_p3[2:0];
  assign xor_ln116_1_fu_1199_p2 = (working_key[4660] == 1'b1)? trunc_ln116_1_fu_1185_p3 ^ select_ln116_1_fu_1173_p3 : trunc_ln116_1_fu_1185_p3 | select_ln116_1_fu_1173_p3;
  assign xor_ln116_fu_1193_p2 = (working_key[4661] == 1'b1)? select_ln116_fu_1165_p3 ^ a_assign_1_fu_1143_p3 : select_ln116_fu_1165_p3 | a_assign_1_fu_1143_p3;
  assign Const_1112 = (1'd1 ^ working_key[4662]);
  assign xor_ln118_1_fu_2281_p2 = (working_key[4663] == 1'b1)? icmp_ln118_1_fu_2107_p2 ^ Const_1112 : icmp_ln118_1_fu_2107_p2 & Const_1112;
  assign Const_1113 = (1'd1 ^ working_key[4664]);
  assign xor_ln118_fu_1377_p2 = (working_key[4665] == 1'b1)? icmp_ln118_reg_4631 ^ Const_1113 : icmp_ln118_reg_4631 << Const_1113;
  assign Const_1114 = (1'd1 ^ working_key[4666]);
  assign xor_ln123_1_fu_2275_p2 = (working_key[4667] == 1'b1)? icmp_ln123_3_fu_2203_p2 ^ Const_1114 : icmp_ln123_3_fu_2203_p2 | Const_1114;
  assign Const_1115 = (1'd1 ^ working_key[4668]);
  assign xor_ln123_fu_1372_p2 = (working_key[4669] == 1'b1)? icmp_ln123_reg_4642 ^ Const_1115 : icmp_ln123_reg_4642 & Const_1115;
  assign Const_1116 = (1'd0 ^ working_key[4670]);
  assign xor_ln155_fu_2619_p2 = (working_key[4671] == 1'b1)? icmp_ln155_fu_2601_p2 << Const_1116 : icmp_ln155_fu_2601_p2 ^ Const_1116;
  assign Const_1117 = (1'd0 ^ working_key[4672]);
  assign xor_ln259_fu_3125_p2 = (working_key[4673] == 1'b1)? icmp_ln259_fu_3073_p2 & Const_1117 : icmp_ln259_fu_3073_p2 ^ Const_1117;
  assign xor_ln95_1_fu_2175_p2 = (working_key[4674] == 1'b1)? trunc_ln116_4_fu_2153_p1 ^ select_ln116_4_fu_2145_p3 : trunc_ln116_4_fu_2153_p1 & select_ln116_4_fu_2145_p3;
  assign xor_ln95_2_fu_2181_p2 = (working_key[4675] == 1'b1)? trunc_ln116_2_fu_2129_p1 & select_ln116_2_fu_2121_p3 : trunc_ln116_2_fu_2129_p1 ^ select_ln116_2_fu_2121_p3;
  assign xor_ln95_3_fu_2187_p2 = (working_key[4676] == 1'b1)? trunc_ln116_3_fu_2141_p1 >> select_ln116_3_fu_2133_p3 : trunc_ln116_3_fu_2141_p1 ^ select_ln116_3_fu_2133_p3;
  assign xor_ln95_fu_2169_p2 = (working_key[4677] == 1'b1)? trunc_ln116_5_fu_2165_p1 ^ select_ln116_5_fu_2157_p3 : trunc_ln116_5_fu_2165_p1 << select_ln116_5_fu_2157_p3;
  assign zext_ln118_fu_2428_p1 = select_ln118_2_fu_2421_p3;
  assign zext_ln123_10_fu_2270_p1 = trunc_ln123_5_fu_2260_p4;
  assign zext_ln123_1_fu_1256_p1 = trunc_ln123_1_fu_1246_p4;
  assign zext_ln123_2_fu_1358_p1 = add_ln123_fu_1352_p2;
  assign zext_ln123_3_fu_1271_p1 = trunc_ln123_2_fu_1261_p4;
  assign zext_ln123_4_fu_2225_p1 = xor_ln95_fu_2169_p2;
  assign zext_ln123_5_fu_2367_p1 = bitoff_q0;
  assign zext_ln123_6_fu_2240_p1 = trunc_ln123_3_fu_2230_p4;
  assign zext_ln123_7_fu_2377_p1 = bitoff_q1;
  assign zext_ln123_8_fu_2255_p1 = trunc_ln123_4_fu_2245_p4;
  assign zext_ln123_9_fu_2393_p1 = add_ln123_4_fu_2387_p2;
  assign zext_ln123_fu_1348_p1 = bitoff_q0;
  assign zext_ln138_1_fu_1866_p1 = add_ln138_1_fu_1860_p2;
  assign zext_ln138_fu_1964_p1 = add_ln138_reg_5073;
  assign zext_ln142_fu_1877_p1 = add_ln142_fu_1871_p2;
  assign zext_ln143_fu_1900_p1 = add_ln143_fu_1894_p2;
  assign zext_ln144_fu_1911_p1 = add_ln144_fu_1905_p2;
  assign zext_ln145_fu_1948_p1 = add_ln145_fu_1942_p2;
  assign zext_ln146_fu_1959_p1 = add_ln146_fu_1953_p2;
  assign zext_ln152_fu_2060_p1 = sext_ln151_fu_2048_p1;
  assign zext_ln187_fu_2455_p1 = i_1_i_reg_928;
  assign zext_ln193_fu_2486_p1 = i_2_i_reg_939;
  assign zext_ln195_fu_2509_p1 = i_3_i_reg_950;
  assign zext_ln206_1_fu_2579_p1 = p_1_rec_i_reg_985;
  assign zext_ln206_fu_2514_p1 = p_1_rec_i_reg_985;
  assign zext_ln225_fu_2793_p1 = m_0_i_reg_1060;
  assign zext_ln226_fu_2804_p1 = m_fu_2798_p2;
  assign zext_ln60_fu_1138_p1 = k_0_i_reg_851;
  assign zext_ln72_fu_2551_p1 = select_ln72_1_fu_2543_p3;
  assign zext_ln75_fu_1520_p1 = lshr_ln76_fu_1514_p2;
  assign zext_ln76_1_fu_1536_p1 = k_1_i_reg_862;
  assign zext_ln76_fu_1510_p1 = add_ln76_fu_1505_p2;
  assign zext_ln89_fu_1566_p1 = sext_ln88_fu_1554_p1;

  always @(posedge ap_clk) begin
    zext_ln75_reg_4696[30:15] <= 16'b0000000000000000;
    sp_0_rec_i_cast_reg_5060[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    zext_ln187_reg_5305[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    zext_ln193_reg_5318[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    zext_ln195_reg_5341[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    zext_ln206_1_reg_5411[4] <= 1'b0;
    zext_ln225_reg_5476[63:32] <= 32'b00000000000000000000000000000000;
  end

  assign working_key = { locking_key[4656:0] };

endmodule



module AddRoundKey_InversMi
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  statemt_address0,
  statemt_ce0,
  statemt_we0,
  statemt_d0,
  statemt_q0,
  statemt_address1,
  statemt_ce1,
  statemt_we1,
  statemt_d1,
  statemt_q1,
  n,
  word_address0,
  word_ce0,
  word_q0,
  word_address1,
  word_ce1,
  word_q1,
  working_key
);

  parameter ap_ST_fsm_state1 = 14'd1;
  parameter ap_ST_fsm_state2 = 14'd2;
  parameter ap_ST_fsm_state3 = 14'd4;
  parameter ap_ST_fsm_state4 = 14'd8;
  parameter ap_ST_fsm_state5 = 14'd16;
  parameter ap_ST_fsm_state6 = 14'd32;
  parameter ap_ST_fsm_state7 = 14'd64;
  parameter ap_ST_fsm_state8 = 14'd128;
  parameter ap_ST_fsm_state9 = 14'd256;
  parameter ap_ST_fsm_state10 = 14'd512;
  parameter ap_ST_fsm_state11 = 14'd1024;
  parameter ap_ST_fsm_state12 = 14'd2048;
  parameter ap_ST_fsm_state13 = 14'd4096;
  parameter ap_ST_fsm_state14 = 14'd8192;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [4:0] statemt_address0;
  output statemt_ce0;
  output statemt_we0;
  output [31:0] statemt_d0;
  input [31:0] statemt_q0;
  output [4:0] statemt_address1;
  output statemt_ce1;
  output statemt_we1;
  output [31:0] statemt_d1;
  input [31:0] statemt_q1;
  input [3:0] n;
  output [8:0] word_address0;
  output word_ce0;
  input [31:0] word_q0;
  output [8:0] word_address1;
  output word_ce1;
  input [31:0] word_q1;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [4:0] statemt_address0;
  reg statemt_ce0;
  reg statemt_we0;
  reg [31:0] statemt_d0;
  reg [4:0] statemt_address1;
  reg statemt_ce1;
  reg statemt_we1;
  reg [31:0] statemt_d1;
  reg [8:0] word_address0;
  reg word_ce0;
  reg [8:0] word_address1;
  reg word_ce1;
  reg [13:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  wire [31:0] grp_fu_320_p2;
  reg [31:0] reg_352;
  wire ap_CS_fsm_state3;
  wire ap_CS_fsm_state4;
  wire [31:0] grp_fu_326_p2;
  reg [31:0] reg_357;
  wire [5:0] tmp_fu_362_p3;
  reg [5:0] tmp_reg_1262;
  wire [2:0] j_2_fu_380_p2;
  reg [2:0] j_2_reg_1270;
  wire ap_CS_fsm_state2;
  wire [5:0] tmp_s_fu_386_p2;
  reg [5:0] tmp_s_reg_1275;
  wire [0:0] exitcond3_fu_374_p2;
  wire [3:0] tmp_4_fu_415_p3;
  reg [3:0] tmp_4_reg_1290;
  reg [4:0] statemt_addr_reg_1296;
  reg [4:0] statemt_addr_17_reg_1301;
  reg [4:0] statemt_addr_18_reg_1316;
  reg [4:0] statemt_addr_19_reg_1321;
  wire [2:0] j_3_fu_490_p2;
  reg [2:0] j_3_reg_1329;
  wire ap_CS_fsm_state6;
  wire [1:0] tmp_2_fu_496_p1;
  reg [1:0] tmp_2_reg_1334;
  wire [0:0] exitcond2_fu_484_p2;
  wire [3:0] tmp_19_fu_500_p3;
  reg [3:0] tmp_19_reg_1341;
  wire [2:0] i_7_fu_518_p2;
  reg [2:0] i_7_reg_1349;
  wire ap_CS_fsm_state7;
  wire [63:0] tmp_30_fu_529_p1;
  reg [63:0] tmp_30_reg_1354;
  wire [0:0] exitcond_fu_512_p2;
  wire [1:0] tmp_45_fu_534_p1;
  reg [1:0] tmp_45_reg_1364;
  wire [30:0] tmp_37_fu_596_p1;
  reg [30:0] tmp_37_reg_1375;
  wire ap_CS_fsm_state8;
  wire [30:0] x_s_fu_600_p2;
  reg [30:0] x_s_reg_1380;
  reg [23:0] tmp_38_reg_1385;
  reg [31:0] statemt_load_20_reg_1390;
  wire [30:0] tmp_56_fu_660_p3;
  reg [30:0] tmp_56_reg_1396;
  reg [23:0] tmp_57_reg_1401;
  reg [31:0] statemt_load_21_reg_1416;
  wire ap_CS_fsm_state9;
  wire [30:0] x_7_fu_926_p2;
  reg [30:0] x_7_reg_1421;
  reg [23:0] tmp_73_reg_1427;
  reg [31:0] statemt_load_22_reg_1432;
  wire [30:0] tmp_90_fu_986_p3;
  reg [30:0] tmp_90_reg_1437;
  reg [23:0] tmp_91_reg_1443;
  wire [31:0] tmp4_fu_1004_p2;
  reg [31:0] tmp4_reg_1448;
  wire [31:0] tmp5_fu_1176_p2;
  reg [31:0] tmp5_reg_1453;
  wire ap_CS_fsm_state10;
  wire [2:0] i_6_fu_1208_p2;
  reg [2:0] i_6_reg_1461;
  wire ap_CS_fsm_state12;
  wire [3:0] tmp_21_fu_1218_p3;
  reg [3:0] tmp_21_reg_1466;
  wire [0:0] exitcond1_fu_1202_p2;
  wire [63:0] tmp_22_fu_1226_p1;
  reg [63:0] tmp_22_reg_1472;
  wire [63:0] tmp_24_fu_1237_p1;
  reg [63:0] tmp_24_reg_1482;
  wire [63:0] tmp_26_fu_1247_p1;
  reg [63:0] tmp_26_reg_1492;
  wire ap_CS_fsm_state13;
  wire [63:0] tmp_28_fu_1257_p1;
  reg [63:0] tmp_28_reg_1502;
  reg [4:0] ret_address0;
  reg ret_ce0;
  reg ret_we0;
  wire [31:0] ret_d0;
  wire [31:0] ret_q0;
  reg [4:0] ret_address1;
  reg ret_ce1;
  wire [31:0] ret_q1;
  reg [2:0] j_reg_276;
  wire ap_CS_fsm_state5;
  reg [2:0] j_1_reg_287;
  reg [2:0] i_reg_298;
  wire ap_CS_fsm_state11;
  reg [2:0] i_1_reg_309;
  wire ap_CS_fsm_state14;
  wire [63:0] tmp_3_fu_391_p1;
  wire [63:0] tmp_16_cast_fu_406_p1;
  wire [63:0] tmp_5_fu_423_p1;
  wire [63:0] tmp_8_fu_434_p1;
  wire [63:0] tmp_17_cast_fu_448_p1;
  wire [63:0] tmp_18_cast_fu_459_p1;
  wire [63:0] tmp_11_fu_469_p1;
  wire [63:0] tmp_14_fu_479_p1;
  wire [63:0] tmp_47_fu_551_p1;
  wire [63:0] tmp_65_fu_690_p1;
  wire [63:0] tmp_82_fu_707_p1;
  wire [5:0] j_cast6_fu_370_p1;
  wire [7:0] tmp_3_cast_fu_396_p1;
  wire [7:0] tmp_16_fu_400_p2;
  wire [1:0] tmp_1_fu_411_p1;
  wire [3:0] tmp_7_fu_428_p2;
  wire [8:0] tmp_3_cast1_fu_439_p1;
  wire [8:0] tmp_17_fu_442_p2;
  wire [8:0] tmp_18_fu_453_p2;
  wire [3:0] tmp_10_fu_464_p2;
  wire [3:0] tmp_13_fu_474_p2;
  wire [3:0] i_cast_fu_508_p1;
  wire [3:0] tmp_29_fu_524_p2;
  wire [1:0] i_7_cast_fu_538_p2;
  wire [3:0] tmp_46_fu_544_p3;
  wire [23:0] grp_fu_332_p4;
  wire [31:0] p_mask_fu_556_p3;
  wire [29:0] tmp_33_fu_570_p1;
  wire [30:0] tmp_34_fu_574_p3;
  wire [0:0] tmp_32_fu_564_p2;
  wire [30:0] tmp_35_fu_582_p2;
  wire [30:0] tmp_36_fu_588_p3;
  wire [23:0] grp_fu_342_p4;
  wire [31:0] p_mask3_fu_616_p3;
  wire [29:0] tmp_51_fu_630_p1;
  wire [30:0] tmp_52_fu_634_p3;
  wire [29:0] tmp_54_fu_648_p1;
  wire [0:0] tmp_50_fu_624_p2;
  wire [30:0] tmp_53_fu_642_p2;
  wire [30:0] tmp_55_fu_652_p3;
  wire [1:0] tmp_97_cast_fu_678_p2;
  wire [3:0] tmp_64_fu_683_p3;
  wire [1:0] tmp_105_cast_fu_695_p2;
  wire [3:0] tmp_81_fu_700_p3;
  wire [31:0] p_mask1_fu_712_p3;
  wire [30:0] tmp_40_fu_725_p2;
  wire [0:0] tmp_39_fu_719_p2;
  wire [30:0] tmp_41_fu_730_p2;
  wire [30:0] tmp_42_fu_736_p3;
  wire [30:0] x_6_fu_744_p2;
  wire [23:0] tmp_43_fu_757_p4;
  wire [31:0] p_mask2_fu_767_p3;
  wire [31:0] x_fu_749_p3;
  wire [0:0] tmp_44_fu_775_p2;
  wire [31:0] x_1_fu_781_p2;
  wire [31:0] p_mask4_fu_798_p3;
  wire [30:0] tmp_59_fu_811_p2;
  wire [0:0] tmp_58_fu_805_p2;
  wire [30:0] tmp_60_fu_816_p2;
  wire [30:0] tmp_61_fu_822_p3;
  wire [30:0] tmp_48_fu_795_p1;
  wire [30:0] x_8_fu_830_p2;
  wire [23:0] tmp_62_fu_844_p4;
  wire [31:0] p_mask5_fu_854_p3;
  wire [31:0] x_3_fu_836_p3;
  wire [0:0] tmp_63_fu_862_p2;
  wire [31:0] x_4_fu_868_p2;
  wire [31:0] p_mask6_fu_882_p3;
  wire [29:0] tmp_68_fu_896_p1;
  wire [30:0] tmp_69_fu_900_p3;
  wire [0:0] tmp_67_fu_890_p2;
  wire [30:0] tmp_70_fu_908_p2;
  wire [30:0] tmp_71_fu_914_p3;
  wire [30:0] tmp_72_fu_922_p1;
  wire [31:0] p_mask9_fu_942_p3;
  wire [29:0] tmp_85_fu_956_p1;
  wire [30:0] tmp_86_fu_960_p3;
  wire [29:0] tmp_88_fu_974_p1;
  wire [0:0] tmp_84_fu_950_p2;
  wire [30:0] tmp_87_fu_968_p2;
  wire [30:0] tmp_89_fu_978_p3;
  wire [31:0] x_2_fu_787_p3;
  wire [31:0] x_5_fu_874_p3;
  wire [31:0] p_mask7_fu_1010_p3;
  wire [30:0] tmp_75_fu_1023_p2;
  wire [0:0] tmp_74_fu_1017_p2;
  wire [30:0] tmp_76_fu_1028_p2;
  wire [30:0] tmp_77_fu_1034_p2;
  wire [30:0] tmp_78_fu_1039_p3;
  wire [23:0] tmp_79_fu_1055_p4;
  wire [31:0] p_mask8_fu_1065_p3;
  wire [31:0] x_9_fu_1047_p3;
  wire [0:0] tmp_80_fu_1073_p2;
  wire [31:0] x_10_fu_1079_p2;
  wire [31:0] p_mask10_fu_1093_p3;
  wire [30:0] tmp_93_fu_1106_p2;
  wire [0:0] tmp_92_fu_1100_p2;
  wire [30:0] tmp_94_fu_1111_p2;
  wire [30:0] tmp_95_fu_1117_p2;
  wire [30:0] tmp_96_fu_1122_p3;
  wire [23:0] tmp_97_fu_1138_p4;
  wire [31:0] p_mask11_fu_1148_p3;
  wire [31:0] x_12_fu_1130_p3;
  wire [0:0] tmp_98_fu_1156_p2;
  wire [31:0] x_13_fu_1162_p2;
  wire [31:0] p_1_fu_1085_p3;
  wire [31:0] x_11_fu_1168_p3;
  wire [31:0] tmp2_fu_1182_p2;
  wire [31:0] tmp3_fu_1191_p2;
  wire [31:0] tmp1_fu_1186_p2;
  wire [1:0] tmp_20_fu_1214_p1;
  wire [3:0] tmp_23_fu_1231_p2;
  wire [3:0] tmp_25_fu_1242_p2;
  wire [3:0] tmp_27_fu_1252_p2;
  reg [13:0] ap_NS_fsm;
  wire [30:0] Const_0;
  wire [30:0] Const_1;
  wire [30:0] Const_2;
  wire [30:0] Const_3;
  wire [30:0] Const_4;
  wire [30:0] Const_5;
  wire [31:0] temp116;
  wire [31:0] temp118;
  wire [31:0] temp119;
  wire [31:0] temp120;
  wire [31:0] temp122;
  wire [31:0] temp123;
  input [12286:0] locking_key;
  wire [209:0] working_key;

  initial begin
    #0 ap_CS_fsm = 14'd1;
  end


  AddRoundKey_Invercud
  #(
    .DataWidth(32),
    .AddressRange(32),
    .AddressWidth(5)
  )
  ret_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(ret_address0),
    .ce0(ret_ce0),
    .we0(ret_we0),
    .d0(ret_d0),
    .q0(ret_q0),
    .address1(ret_address1),
    .ce1(ret_ce1),
    .q1(ret_q1)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state6) & (exitcond2_fu_484_p2 == 1'd1)) begin
      if(working_key[200] == 1'b1) begin
        i_1_reg_309 <= temp116;
      end else begin
        i_1_reg_309 <= 3'd0;
      end
    end else if(1'b1 == ap_CS_fsm_state14) begin
      i_1_reg_309 <= i_6_reg_1461;
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond2_fu_484_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state6)) begin
      if(working_key[203] == 1'b1) begin
        i_reg_298 <= 3'd0;
      end else begin
        i_reg_298 <= temp120;
      end
    end else if(1'b1 == ap_CS_fsm_state11) begin
      i_reg_298 <= i_7_reg_1349;
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond3_fu_374_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
      j_1_reg_287 <= 3'd0;
    end else if((1'b1 == ap_CS_fsm_state7) & (exitcond_fu_512_p2 == 1'd1)) begin
      j_1_reg_287 <= j_3_reg_1329;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      j_reg_276 <= j_2_reg_1270;
    end else if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      j_reg_276 <= 3'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      i_6_reg_1461 <= i_6_fu_1208_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      i_7_reg_1349 <= i_7_fu_518_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      j_2_reg_1270 <= j_2_fu_380_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state6) begin
      j_3_reg_1329 <= j_3_fu_490_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3)) begin
      reg_352 <= grp_fu_320_p2;
      reg_357 <= grp_fu_326_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond3_fu_374_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      statemt_addr_17_reg_1301[3:2] <= tmp_8_fu_434_p1[3:2];
      statemt_addr_reg_1296[3:2] <= tmp_5_fu_423_p1[3:2];
      tmp_4_reg_1290[3:2] <= tmp_4_fu_415_p3[3:2];
      tmp_s_reg_1275 <= tmp_s_fu_386_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      statemt_addr_18_reg_1316[3:2] <= tmp_11_fu_469_p1[3:2];
      statemt_addr_19_reg_1321[3:2] <= tmp_14_fu_479_p1[3:2];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state8) begin
      statemt_load_20_reg_1390 <= statemt_q1;
      tmp_37_reg_1375 <= tmp_37_fu_596_p1;
      tmp_38_reg_1385 <= { { x_s_fu_600_p2[30:7] } };
      tmp_56_reg_1396 <= tmp_56_fu_660_p3;
      tmp_57_reg_1401 <= { { tmp_56_fu_660_p3[30:7] } };
      x_s_reg_1380 <= x_s_fu_600_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      statemt_load_21_reg_1416 <= statemt_q0;
      statemt_load_22_reg_1432 <= statemt_q1;
      tmp4_reg_1448 <= tmp4_fu_1004_p2;
      tmp_73_reg_1427 <= { { x_7_fu_926_p2[30:7] } };
      tmp_90_reg_1437 <= tmp_90_fu_986_p3;
      tmp_91_reg_1443 <= { { tmp_90_fu_986_p3[30:7] } };
      x_7_reg_1421 <= x_7_fu_926_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state10) begin
      tmp5_reg_1453 <= tmp5_fu_1176_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond2_fu_484_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state6)) begin
      tmp_19_reg_1341[3:2] <= tmp_19_fu_500_p3[3:2];
      tmp_2_reg_1334 <= tmp_2_fu_496_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond1_fu_1202_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state12)) begin
      tmp_21_reg_1466[3:2] <= tmp_21_fu_1218_p3[3:2];
      tmp_22_reg_1472[3:2] <= tmp_22_fu_1226_p1[3:2];
      tmp_24_reg_1482[3:2] <= tmp_24_fu_1237_p1[3:2];
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      tmp_26_reg_1492[3:2] <= tmp_26_fu_1247_p1[3:2];
      tmp_28_reg_1502[3:2] <= tmp_28_fu_1257_p1[3:2];
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond_fu_512_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      tmp_30_reg_1354[3:0] <= tmp_30_fu_529_p1[3:0];
      tmp_45_reg_1364 <= tmp_45_fu_534_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      tmp_reg_1262[5:2] <= tmp_fu_362_p3[5:2];
    end 
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1) | (1'b1 == ap_CS_fsm_state12) & (exitcond1_fu_1202_p2 == 1'd1)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state12) & (exitcond1_fu_1202_p2 == 1'd1)) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      ret_address0 = tmp_28_fu_1257_p1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      ret_address0 = tmp_22_fu_1226_p1;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      ret_address0 = tmp_30_reg_1354;
    end else begin
      ret_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      ret_address1 = tmp_26_fu_1247_p1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      ret_address1 = tmp_24_fu_1237_p1;
    end else begin
      ret_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12)) begin
      ret_ce0 = 1'b1;
    end else begin
      ret_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12)) begin
      ret_ce1 = 1'b1;
    end else begin
      ret_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      ret_we0 = 1'b1;
    end else begin
      ret_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state14) begin
      statemt_address0 = tmp_26_reg_1492;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_address0 = tmp_22_reg_1472;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address0 = tmp_65_fu_690_p1;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      statemt_address0 = tmp_30_fu_529_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address0 = statemt_addr_18_reg_1316;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address0 = statemt_addr_reg_1296;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address0 = tmp_11_fu_469_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address0 = tmp_5_fu_423_p1;
    end else begin
      statemt_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state14) begin
      statemt_address1 = tmp_28_reg_1502;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_address1 = tmp_24_reg_1482;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address1 = tmp_82_fu_707_p1;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      statemt_address1 = tmp_47_fu_551_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address1 = statemt_addr_19_reg_1321;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address1 = statemt_addr_17_reg_1301;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address1 = tmp_14_fu_479_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address1 = tmp_8_fu_434_p1;
    end else begin
      statemt_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7)) begin
      statemt_ce0 = 1'b1;
    end else begin
      statemt_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7)) begin
      statemt_ce1 = 1'b1;
    end else begin
      statemt_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state14) begin
      statemt_d0 = ret_q1;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_d0 = ret_q0;
    end else if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5)) begin
      statemt_d0 = reg_352;
    end else begin
      statemt_d0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state14) begin
      statemt_d1 = ret_q0;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_d1 = ret_q1;
    end else if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5)) begin
      statemt_d1 = reg_357;
    end else begin
      statemt_d1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state13)) begin
      statemt_we0 = 1'b1;
    end else begin
      statemt_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state13)) begin
      statemt_we1 = 1'b1;
    end else begin
      statemt_we1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      word_address0 = tmp_17_cast_fu_448_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      word_address0 = tmp_3_fu_391_p1;
    end else begin
      word_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      word_address1 = tmp_18_cast_fu_459_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      word_address1 = tmp_16_cast_fu_406_p1;
    end else begin
      word_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state3)) begin
      word_ce0 = 1'b1;
    end else begin
      word_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state3)) begin
      word_ce1 = 1'b1;
    end else begin
      word_ce1 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if((exitcond3_fu_374_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end
      end
      ap_ST_fsm_state3: begin
        ap_NS_fsm = ap_ST_fsm_state4;
      end
      ap_ST_fsm_state4: begin
        ap_NS_fsm = ap_ST_fsm_state5;
      end
      ap_ST_fsm_state5: begin
        ap_NS_fsm = ap_ST_fsm_state2;
      end
      ap_ST_fsm_state6: begin
        if((1'b1 == ap_CS_fsm_state6) & (exitcond2_fu_484_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state12;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end
      end
      ap_ST_fsm_state7: begin
        if((1'b1 == ap_CS_fsm_state7) & (exitcond_fu_512_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state8: begin
        ap_NS_fsm = ap_ST_fsm_state9;
      end
      ap_ST_fsm_state9: begin
        ap_NS_fsm = ap_ST_fsm_state10;
      end
      ap_ST_fsm_state10: begin
        ap_NS_fsm = ap_ST_fsm_state11;
      end
      ap_ST_fsm_state11: begin
        ap_NS_fsm = ap_ST_fsm_state7;
      end
      ap_ST_fsm_state12: begin
        if((1'b1 == ap_CS_fsm_state12) & (exitcond1_fu_1202_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state13;
        end
      end
      ap_ST_fsm_state13: begin
        ap_NS_fsm = ap_ST_fsm_state14;
      end
      ap_ST_fsm_state14: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign exitcond1_fu_1202_p2 = (i_1_reg_309 == 3'd4)? 1'b1 : 1'b0;
  assign exitcond2_fu_484_p2 = (j_1_reg_287 == 3'd4)? 1'b1 : 1'b0;
  assign exitcond3_fu_374_p2 = (j_reg_276 == 3'd4)? 1'b1 : 1'b0;
  assign exitcond_fu_512_p2 = (i_reg_298 == 3'd4)? 1'b1 : 1'b0;
  assign grp_fu_320_p2 = word_q0 ^ statemt_q0;
  assign grp_fu_326_p2 = word_q1 ^ statemt_q1;
  assign grp_fu_332_p4 = { { statemt_q0[30:7] } };
  assign grp_fu_342_p4 = { { statemt_q1[30:7] } };
  assign i_6_fu_1208_p2 = i_1_reg_309 + 3'd1;
  assign i_7_cast_fu_538_p2 = tmp_45_fu_534_p1 + 2'd1;
  assign i_7_fu_518_p2 = i_reg_298 + 3'd1;
  assign i_cast_fu_508_p1 = i_reg_298;
  assign j_2_fu_380_p2 = j_reg_276 + 3'd1;
  assign j_3_fu_490_p2 = j_1_reg_287 + 3'd1;
  assign j_cast6_fu_370_p1 = j_reg_276;
  assign p_1_fu_1085_p3 = (tmp_80_fu_1073_p2[0:0] === 1'b1)? x_10_fu_1079_p2 : x_9_fu_1047_p3;
  assign p_mask10_fu_1093_p3 = { { tmp_91_reg_1443 }, { 8'd0 } };
  assign p_mask11_fu_1148_p3 = { { tmp_97_fu_1138_p4 }, { 8'd0 } };
  assign p_mask1_fu_712_p3 = { { tmp_38_reg_1385 }, { 8'd0 } };
  assign p_mask2_fu_767_p3 = { { tmp_43_fu_757_p4 }, { 8'd0 } };
  assign p_mask3_fu_616_p3 = { { grp_fu_342_p4 }, { 8'd0 } };
  assign p_mask4_fu_798_p3 = { { tmp_57_reg_1401 }, { 8'd0 } };
  assign p_mask5_fu_854_p3 = { { tmp_62_fu_844_p4 }, { 8'd0 } };
  assign p_mask6_fu_882_p3 = { { grp_fu_332_p4 }, { 8'd0 } };
  assign p_mask7_fu_1010_p3 = { { tmp_73_reg_1427 }, { 8'd0 } };
  assign p_mask8_fu_1065_p3 = { { tmp_79_fu_1055_p4 }, { 8'd0 } };
  assign p_mask9_fu_942_p3 = { { grp_fu_342_p4 }, { 8'd0 } };
  assign p_mask_fu_556_p3 = { { grp_fu_332_p4 }, { 8'd0 } };
  assign ret_d0 = tmp3_fu_1191_p2 ^ tmp1_fu_1186_p2;
  assign tmp1_fu_1186_p2 = tmp2_fu_1182_p2 ^ statemt_load_20_reg_1390;
  assign tmp2_fu_1182_p2 = statemt_load_22_reg_1432 ^ statemt_load_21_reg_1416;
  assign tmp3_fu_1191_p2 = tmp5_reg_1453 ^ tmp4_reg_1448;
  assign tmp4_fu_1004_p2 = x_5_fu_874_p3 ^ x_2_fu_787_p3;
  assign tmp5_fu_1176_p2 = x_11_fu_1168_p3 ^ p_1_fu_1085_p3;
  assign tmp_105_cast_fu_695_p2 = $signed(tmp_45_reg_1364) + $signed(2'd3);
  assign tmp_10_fu_464_p2 = tmp_4_reg_1290 | 4'd2;
  assign tmp_11_fu_469_p1 = tmp_10_fu_464_p2;
  assign tmp_13_fu_474_p2 = tmp_4_reg_1290 | 4'd3;
  assign tmp_14_fu_479_p1 = tmp_13_fu_474_p2;
  assign tmp_16_cast_fu_406_p1 = tmp_16_fu_400_p2;
  assign tmp_16_fu_400_p2 = 8'd120 + tmp_3_cast_fu_396_p1;
  assign tmp_17_cast_fu_448_p1 = tmp_17_fu_442_p2;
  assign tmp_17_fu_442_p2 = 9'd240 + tmp_3_cast1_fu_439_p1;
  assign tmp_18_cast_fu_459_p1 = tmp_18_fu_453_p2;
  assign tmp_18_fu_453_p2 = $signed(9'd360) + $signed(tmp_3_cast1_fu_439_p1);
  assign tmp_19_fu_500_p3 = { { tmp_2_fu_496_p1 }, { 2'd0 } };
  assign tmp_1_fu_411_p1 = j_reg_276[1:0];
  assign tmp_20_fu_1214_p1 = i_1_reg_309[1:0];
  assign tmp_21_fu_1218_p3 = { { tmp_20_fu_1214_p1 }, { 2'd0 } };
  assign tmp_22_fu_1226_p1 = tmp_21_fu_1218_p3;
  assign tmp_23_fu_1231_p2 = tmp_21_fu_1218_p3 | 4'd1;
  assign tmp_24_fu_1237_p1 = tmp_23_fu_1231_p2;
  assign tmp_25_fu_1242_p2 = tmp_21_reg_1466 | 4'd2;
  assign tmp_26_fu_1247_p1 = tmp_25_fu_1242_p2;
  assign tmp_27_fu_1252_p2 = tmp_21_reg_1466 | 4'd3;
  assign tmp_28_fu_1257_p1 = tmp_27_fu_1252_p2;
  assign tmp_29_fu_524_p2 = tmp_19_reg_1341 + i_cast_fu_508_p1;
  assign tmp_2_fu_496_p1 = j_1_reg_287[1:0];
  assign tmp_30_fu_529_p1 = tmp_29_fu_524_p2;
  assign tmp_32_fu_564_p2 = (p_mask_fu_556_p3 == 32'd256)? 1'b1 : 1'b0;
  assign tmp_33_fu_570_p1 = statemt_q0[29:0];
  assign tmp_34_fu_574_p3 = { { tmp_33_fu_570_p1 }, { 1'd0 } };
  assign tmp_35_fu_582_p2 = tmp_34_fu_574_p3 ^ 31'd283;
  assign tmp_36_fu_588_p3 = (tmp_32_fu_564_p2[0:0] === 1'b1)? tmp_35_fu_582_p2 : tmp_34_fu_574_p3;
  assign tmp_37_fu_596_p1 = statemt_q0[30:0];
  assign tmp_39_fu_719_p2 = (p_mask1_fu_712_p3 == 32'd256)? 1'b1 : 1'b0;
  assign tmp_3_cast1_fu_439_p1 = tmp_s_reg_1275;
  assign tmp_3_cast_fu_396_p1 = tmp_s_fu_386_p2;
  assign tmp_3_fu_391_p1 = tmp_s_fu_386_p2;
  assign Const_0 = (31'd1398052267 ^ working_key[42:12]);
  assign tmp_40_fu_725_p2 = x_s_reg_1380 << Const_0;
  assign tmp_41_fu_730_p2 = tmp_40_fu_725_p2 ^ 31'd283;
  assign tmp_42_fu_736_p3 = (tmp_39_fu_719_p2[0:0] === 1'b1)? tmp_41_fu_730_p2 : tmp_40_fu_725_p2;
  assign tmp_43_fu_757_p4 = { { x_6_fu_744_p2[30:7] } };
  assign tmp_44_fu_775_p2 = (p_mask2_fu_767_p3 == 32'd256)? 1'b1 : 1'b0;
  assign tmp_45_fu_534_p1 = i_reg_298[1:0];
  assign tmp_46_fu_544_p3 = { { tmp_2_reg_1334 }, { i_7_cast_fu_538_p2 } };
  assign tmp_47_fu_551_p1 = tmp_46_fu_544_p3;
  assign tmp_48_fu_795_p1 = statemt_load_20_reg_1390[30:0];
  assign tmp_4_fu_415_p3 = { { tmp_1_fu_411_p1 }, { 2'd0 } };
  assign tmp_50_fu_624_p2 = (p_mask3_fu_616_p3 == 32'd256)? 1'b1 : 1'b0;
  assign tmp_51_fu_630_p1 = statemt_q1[29:0];
  assign tmp_52_fu_634_p3 = { { tmp_51_fu_630_p1 }, { 1'd0 } };
  assign tmp_53_fu_642_p2 = tmp_52_fu_634_p3 ^ 31'd283;
  assign tmp_54_fu_648_p1 = statemt_q1[29:0];
  assign tmp_55_fu_652_p3 = { { tmp_54_fu_648_p1 }, { 1'd0 } };
  assign tmp_56_fu_660_p3 = (tmp_50_fu_624_p2[0:0] === 1'b1)? tmp_53_fu_642_p2 : tmp_55_fu_652_p3;
  assign tmp_58_fu_805_p2 = (p_mask4_fu_798_p3 == 32'd256)? 1'b1 : 1'b0;
  assign Const_1 = (31'd1297241770 ^ working_key[73:43]);
  assign tmp_59_fu_811_p2 = tmp_56_reg_1396 << Const_1;
  assign tmp_5_fu_423_p1 = tmp_4_fu_415_p3;
  assign tmp_60_fu_816_p2 = tmp_59_fu_811_p2 ^ 31'd283;
  assign tmp_61_fu_822_p3 = (tmp_58_fu_805_p2[0:0] === 1'b1)? tmp_60_fu_816_p2 : tmp_59_fu_811_p2;
  assign tmp_62_fu_844_p4 = { { x_8_fu_830_p2[30:7] } };
  assign tmp_63_fu_862_p2 = (p_mask5_fu_854_p3 == 32'd256)? 1'b1 : 1'b0;
  assign tmp_64_fu_683_p3 = { { tmp_2_reg_1334 }, { tmp_97_cast_fu_678_p2 } };
  assign tmp_65_fu_690_p1 = tmp_64_fu_683_p3;
  assign tmp_67_fu_890_p2 = (p_mask6_fu_882_p3 == 32'd256)? 1'b1 : 1'b0;
  assign tmp_68_fu_896_p1 = statemt_q0[29:0];
  assign tmp_69_fu_900_p3 = { { tmp_68_fu_896_p1 }, { 1'd0 } };
  assign tmp_70_fu_908_p2 = tmp_69_fu_900_p3 ^ 31'd283;
  assign tmp_71_fu_914_p3 = (tmp_67_fu_890_p2[0:0] === 1'b1)? tmp_70_fu_908_p2 : tmp_69_fu_900_p3;
  assign tmp_72_fu_922_p1 = statemt_q0[30:0];
  assign tmp_74_fu_1017_p2 = (p_mask7_fu_1010_p3 == 32'd256)? 1'b1 : 1'b0;
  assign Const_2 = (31'd1431644927 ^ working_key[104:74]);
  assign tmp_75_fu_1023_p2 = x_7_reg_1421 << Const_2;
  assign tmp_76_fu_1028_p2 = tmp_75_fu_1023_p2 ^ 31'd283;
  assign Const_3 = (31'd715827723 ^ working_key[135:105]);
  assign tmp_77_fu_1034_p2 = x_7_reg_1421 << Const_3;
  assign tmp_78_fu_1039_p3 = (tmp_74_fu_1017_p2[0:0] === 1'b1)? tmp_76_fu_1028_p2 : tmp_77_fu_1034_p2;
  assign tmp_79_fu_1055_p4 = { { tmp_78_fu_1039_p3[30:7] } };
  assign tmp_7_fu_428_p2 = tmp_4_fu_415_p3 | 4'd1;
  assign tmp_80_fu_1073_p2 = (p_mask8_fu_1065_p3 == 32'd256)? 1'b1 : 1'b0;
  assign tmp_81_fu_700_p3 = { { tmp_2_reg_1334 }, { tmp_105_cast_fu_695_p2 } };
  assign tmp_82_fu_707_p1 = tmp_81_fu_700_p3;
  assign tmp_84_fu_950_p2 = (p_mask9_fu_942_p3 == 32'd256)? 1'b1 : 1'b0;
  assign tmp_85_fu_956_p1 = statemt_q1[29:0];
  assign tmp_86_fu_960_p3 = { { tmp_85_fu_956_p1 }, { 1'd0 } };
  assign tmp_87_fu_968_p2 = tmp_86_fu_960_p3 ^ 31'd283;
  assign tmp_88_fu_974_p1 = statemt_q1[29:0];
  assign tmp_89_fu_978_p3 = { { tmp_88_fu_974_p1 }, { 1'd0 } };
  assign tmp_8_fu_434_p1 = tmp_7_fu_428_p2;
  assign tmp_90_fu_986_p3 = (tmp_84_fu_950_p2[0:0] === 1'b1)? tmp_87_fu_968_p2 : tmp_89_fu_978_p3;
  assign tmp_92_fu_1100_p2 = (p_mask10_fu_1093_p3 == 32'd256)? 1'b1 : 1'b0;
  assign Const_4 = (31'd893999783 ^ working_key[166:136]);
  assign tmp_93_fu_1106_p2 = tmp_90_reg_1437 << Const_4;
  assign tmp_94_fu_1111_p2 = tmp_93_fu_1106_p2 ^ 31'd283;
  assign Const_5 = (31'd1428515515 ^ working_key[197:167]);
  assign tmp_95_fu_1117_p2 = tmp_90_reg_1437 << Const_5;
  assign tmp_96_fu_1122_p3 = (tmp_92_fu_1100_p2[0:0] === 1'b1)? tmp_94_fu_1111_p2 : tmp_95_fu_1117_p2;
  assign tmp_97_cast_fu_678_p2 = tmp_45_reg_1364 ^ 2'd2;
  assign tmp_97_fu_1138_p4 = { { tmp_96_fu_1122_p3[30:7] } };
  assign tmp_98_fu_1156_p2 = (p_mask11_fu_1148_p3 == 32'd256)? 1'b1 : 1'b0;
  assign tmp_fu_362_p3 = { { n }, { 2'd0 } };
  assign tmp_s_fu_386_p2 = j_cast6_fu_370_p1 + tmp_reg_1262;
  assign x_10_fu_1079_p2 = x_9_fu_1047_p3 ^ 32'd283;
  assign x_11_fu_1168_p3 = (tmp_98_fu_1156_p2[0:0] === 1'b1)? x_13_fu_1162_p2 : x_12_fu_1130_p3;
  assign x_12_fu_1130_p3 = { { tmp_96_fu_1122_p3 }, { 1'd0 } };
  assign x_13_fu_1162_p2 = x_12_fu_1130_p3 ^ 32'd283;
  assign x_1_fu_781_p2 = x_fu_749_p3 ^ 32'd283;
  assign x_2_fu_787_p3 = (tmp_44_fu_775_p2[0:0] === 1'b1)? x_1_fu_781_p2 : x_fu_749_p3;
  assign x_3_fu_836_p3 = { { x_8_fu_830_p2 }, { 1'd0 } };
  assign x_4_fu_868_p2 = x_3_fu_836_p3 ^ 32'd283;
  assign x_5_fu_874_p3 = (tmp_63_fu_862_p2[0:0] === 1'b1)? x_4_fu_868_p2 : x_3_fu_836_p3;
  assign x_6_fu_744_p2 = tmp_42_fu_736_p3 ^ tmp_37_reg_1375;
  assign x_7_fu_926_p2 = tmp_72_fu_922_p1 ^ tmp_71_fu_914_p3;
  assign x_8_fu_830_p2 = tmp_61_fu_822_p3 ^ tmp_48_fu_795_p1;
  assign x_9_fu_1047_p3 = { { tmp_78_fu_1039_p3 }, { 1'd0 } };
  assign x_fu_749_p3 = { { x_6_fu_744_p2 }, { 1'd0 } };
  assign x_s_fu_600_p2 = tmp_37_fu_596_p1 ^ tmp_36_fu_588_p3;

  always @(posedge ap_clk) begin
    tmp_reg_1262[1:0] <= 2'b00;
    tmp_4_reg_1290[1:0] <= 2'b00;
    statemt_addr_reg_1296[1:0] <= 2'b00;
    statemt_addr_reg_1296[4] <= 1'b0;
    statemt_addr_17_reg_1301[1:0] <= 2'b01;
    statemt_addr_17_reg_1301[4] <= 1'b0;
    statemt_addr_18_reg_1316[1:0] <= 2'b10;
    statemt_addr_18_reg_1316[4] <= 1'b0;
    statemt_addr_19_reg_1321[1:0] <= 2'b11;
    statemt_addr_19_reg_1321[4] <= 1'b0;
    tmp_19_reg_1341[1:0] <= 2'b00;
    tmp_30_reg_1354[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    tmp_21_reg_1466[1:0] <= 2'b00;
    tmp_22_reg_1472[1:0] <= 2'b00;
    tmp_22_reg_1472[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    tmp_24_reg_1482[1:0] <= 2'b01;
    tmp_24_reg_1482[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    tmp_26_reg_1492[1:0] <= 2'b10;
    tmp_26_reg_1492[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    tmp_28_reg_1502[1:0] <= 2'b11;
    tmp_28_reg_1502[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
  end

  assign temp116 = temp118 * temp119;
  assign temp119 = (working_key[198] == 1'b1)? statemt_q0 + statemt_q1 : word_q0 + word_q1;
  assign temp118 = (working_key[199] == 1'b1)? statemt_q1 + word_q1 : statemt_q1 + word_q1;
  assign temp120 = temp122 * temp123;
  assign temp123 = (working_key[201] == 1'b1)? word_q0 + statemt_q0 : statemt_q1 + word_q0;
  assign temp122 = (working_key[202] == 1'b1)? n + word_q1 : n + word_q0;
  assign working_key = { locking_key[187:0] };

endmodule



module aes_func_call_en
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  statemt1_address0,
  statemt1_ce0,
  statemt1_we0,
  statemt1_d0,
  statemt1_q0,
  working_key
);

  parameter ap_ST_fsm_state1 = 13'd1;
  parameter ap_ST_fsm_state2 = 13'd2;
  parameter ap_ST_fsm_state3 = 13'd4;
  parameter ap_ST_fsm_state4 = 13'd8;
  parameter ap_ST_fsm_state5 = 13'd16;
  parameter ap_ST_fsm_state6 = 13'd32;
  parameter ap_ST_fsm_state7 = 13'd64;
  parameter ap_ST_fsm_state8 = 13'd128;
  parameter ap_ST_fsm_state9 = 13'd256;
  parameter ap_ST_fsm_state10 = 13'd512;
  parameter ap_ST_fsm_state11 = 13'd1024;
  parameter ap_ST_fsm_state12 = 13'd2048;
  parameter ap_ST_fsm_state13 = 13'd4096;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [4:0] statemt1_address0;
  output statemt1_ce0;
  output statemt1_we0;
  output [31:0] statemt1_d0;
  input [31:0] statemt1_q0;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [4:0] statemt1_address0;
  reg statemt1_ce0;
  reg statemt1_we0;
  reg [12:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  wire [5:0] i_3_fu_154_p2;
  reg [5:0] i_3_reg_197;
  wire ap_CS_fsm_state2;
  wire [63:0] tmp_fu_160_p1;
  reg [63:0] tmp_reg_202;
  wire [0:0] exitcond6_fu_148_p2;
  wire [3:0] i_4_fu_171_p2;
  reg [3:0] i_4_reg_215;
  wire ap_CS_fsm_state7;
  wire [5:0] i_5_fu_183_p2;
  reg [5:0] i_5_reg_223;
  wire ap_CS_fsm_state12;
  wire [63:0] tmp_3_fu_189_p1;
  reg [63:0] tmp_3_reg_228;
  wire [0:0] exitcond_fu_177_p2;
  reg [4:0] statemt_address0;
  reg statemt_ce0;
  reg statemt_we0;
  reg [31:0] statemt_d0;
  wire [31:0] statemt_q0;
  reg [4:0] statemt_address1;
  reg statemt_ce1;
  reg statemt_we1;
  reg [31:0] statemt_d1;
  wire [31:0] statemt_q1;
  wire grp_MixColumn_AddRoundKe_fu_122_ap_start;
  wire grp_MixColumn_AddRoundKe_fu_122_ap_done;
  wire grp_MixColumn_AddRoundKe_fu_122_ap_idle;
  wire grp_MixColumn_AddRoundKe_fu_122_ap_ready;
  wire [4:0] grp_MixColumn_AddRoundKe_fu_122_statemt_address0;
  wire grp_MixColumn_AddRoundKe_fu_122_statemt_ce0;
  wire grp_MixColumn_AddRoundKe_fu_122_statemt_we0;
  wire [31:0] grp_MixColumn_AddRoundKe_fu_122_statemt_d0;
  wire [4:0] grp_MixColumn_AddRoundKe_fu_122_statemt_address1;
  wire grp_MixColumn_AddRoundKe_fu_122_statemt_ce1;
  wire grp_MixColumn_AddRoundKe_fu_122_statemt_we1;
  wire [31:0] grp_MixColumn_AddRoundKe_fu_122_statemt_d1;
  wire grp_ByteSub_ShiftRow_fu_131_ap_start;
  wire grp_ByteSub_ShiftRow_fu_131_ap_done;
  wire grp_ByteSub_ShiftRow_fu_131_ap_idle;
  wire grp_ByteSub_ShiftRow_fu_131_ap_ready;
  wire [4:0] grp_ByteSub_ShiftRow_fu_131_statemt_address0;
  wire grp_ByteSub_ShiftRow_fu_131_statemt_ce0;
  wire grp_ByteSub_ShiftRow_fu_131_statemt_we0;
  wire [31:0] grp_ByteSub_ShiftRow_fu_131_statemt_d0;
  wire [4:0] grp_ByteSub_ShiftRow_fu_131_statemt_address1;
  wire grp_ByteSub_ShiftRow_fu_131_statemt_ce1;
  wire grp_ByteSub_ShiftRow_fu_131_statemt_we1;
  wire [31:0] grp_ByteSub_ShiftRow_fu_131_statemt_d1;
  wire grp_AddRoundKey_fu_138_ap_start;
  wire grp_AddRoundKey_fu_138_ap_done;
  wire grp_AddRoundKey_fu_138_ap_idle;
  wire grp_AddRoundKey_fu_138_ap_ready;
  wire [4:0] grp_AddRoundKey_fu_138_statemt_address0;
  wire grp_AddRoundKey_fu_138_statemt_ce0;
  wire grp_AddRoundKey_fu_138_statemt_we0;
  wire [31:0] grp_AddRoundKey_fu_138_statemt_d0;
  wire [4:0] grp_AddRoundKey_fu_138_statemt_address1;
  wire grp_AddRoundKey_fu_138_statemt_ce1;
  wire grp_AddRoundKey_fu_138_statemt_we1;
  wire [31:0] grp_AddRoundKey_fu_138_statemt_d1;
  reg [5:0] grp_AddRoundKey_fu_138_n;
  reg [5:0] i_reg_88;
  wire ap_CS_fsm_state3;
  reg [3:0] i_1_reg_99;
  wire ap_CS_fsm_state8;
  wire ap_CS_fsm_state4;
  reg [5:0] i_2_reg_111;
  wire ap_CS_fsm_state13;
  wire ap_CS_fsm_state11;
  reg grp_MixColumn_AddRoundKe_fu_122_ap_start_reg;
  reg grp_ByteSub_ShiftRow_fu_131_ap_start_reg;
  wire ap_CS_fsm_state5;
  wire [0:0] exitcond7_fu_165_p2;
  wire ap_CS_fsm_state6;
  wire ap_CS_fsm_state9;
  reg grp_AddRoundKey_fu_138_ap_start_reg;
  wire ap_CS_fsm_state10;
  reg [12:0] ap_NS_fsm;
  wire [31:0] temp100;
  wire [31:0] temp102;
  wire [31:0] temp103;
  wire [31:0] temp104;
  wire [31:0] temp106;
  wire [31:0] temp107;
  input [23:0] working_key;

  initial begin
    #0 ap_CS_fsm = 13'd1;
    #0 grp_MixColumn_AddRoundKe_fu_122_ap_start_reg = 1'b0;
    #0 grp_ByteSub_ShiftRow_fu_131_ap_start_reg = 1'b0;
    #0 grp_AddRoundKey_fu_138_ap_start_reg = 1'b0;
  end


  MixColumn_AddRoundEe
  #(
    .DataWidth(32),
    .AddressRange(32),
    .AddressWidth(5)
  )
  statemt_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(statemt_address0),
    .ce0(statemt_ce0),
    .we0(statemt_we0),
    .d0(statemt_d0),
    .q0(statemt_q0),
    .address1(statemt_address1),
    .ce1(statemt_ce1),
    .we1(statemt_we1),
    .d1(statemt_d1),
    .q1(statemt_q1)
  );


  MixColumn_AddRoundKe
  grp_MixColumn_AddRoundKe_fu_122
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_MixColumn_AddRoundKe_fu_122_ap_start),
    .ap_done(grp_MixColumn_AddRoundKe_fu_122_ap_done),
    .ap_idle(grp_MixColumn_AddRoundKe_fu_122_ap_idle),
    .ap_ready(grp_MixColumn_AddRoundKe_fu_122_ap_ready),
    .statemt_address0(grp_MixColumn_AddRoundKe_fu_122_statemt_address0),
    .statemt_ce0(grp_MixColumn_AddRoundKe_fu_122_statemt_ce0),
    .statemt_we0(grp_MixColumn_AddRoundKe_fu_122_statemt_we0),
    .statemt_d0(grp_MixColumn_AddRoundKe_fu_122_statemt_d0),
    .statemt_q0(statemt_q0),
    .statemt_address1(grp_MixColumn_AddRoundKe_fu_122_statemt_address1),
    .statemt_ce1(grp_MixColumn_AddRoundKe_fu_122_statemt_ce1),
    .statemt_we1(grp_MixColumn_AddRoundKe_fu_122_statemt_we1),
    .statemt_d1(grp_MixColumn_AddRoundKe_fu_122_statemt_d1),
    .statemt_q1(statemt_q1),
    .n(i_1_reg_99),
    .working_key(working_key)
  );


  ByteSub_ShiftRow
  grp_ByteSub_ShiftRow_fu_131
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_ByteSub_ShiftRow_fu_131_ap_start),
    .ap_done(grp_ByteSub_ShiftRow_fu_131_ap_done),
    .ap_idle(grp_ByteSub_ShiftRow_fu_131_ap_idle),
    .ap_ready(grp_ByteSub_ShiftRow_fu_131_ap_ready),
    .statemt_address0(grp_ByteSub_ShiftRow_fu_131_statemt_address0),
    .statemt_ce0(grp_ByteSub_ShiftRow_fu_131_statemt_ce0),
    .statemt_we0(grp_ByteSub_ShiftRow_fu_131_statemt_we0),
    .statemt_d0(grp_ByteSub_ShiftRow_fu_131_statemt_d0),
    .statemt_q0(statemt_q0),
    .statemt_address1(grp_ByteSub_ShiftRow_fu_131_statemt_address1),
    .statemt_ce1(grp_ByteSub_ShiftRow_fu_131_statemt_ce1),
    .statemt_we1(grp_ByteSub_ShiftRow_fu_131_statemt_we1),
    .statemt_d1(grp_ByteSub_ShiftRow_fu_131_statemt_d1),
    .statemt_q1(statemt_q1),
    .working_key(working_key)
  );


  AddRoundKey
  grp_AddRoundKey_fu_138
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_AddRoundKey_fu_138_ap_start),
    .ap_done(grp_AddRoundKey_fu_138_ap_done),
    .ap_idle(grp_AddRoundKey_fu_138_ap_idle),
    .ap_ready(grp_AddRoundKey_fu_138_ap_ready),
    .statemt_address0(grp_AddRoundKey_fu_138_statemt_address0),
    .statemt_ce0(grp_AddRoundKey_fu_138_statemt_ce0),
    .statemt_we0(grp_AddRoundKey_fu_138_statemt_we0),
    .statemt_d0(grp_AddRoundKey_fu_138_statemt_d0),
    .statemt_q0(statemt_q0),
    .statemt_address1(grp_AddRoundKey_fu_138_statemt_address1),
    .statemt_ce1(grp_AddRoundKey_fu_138_statemt_ce1),
    .statemt_we1(grp_AddRoundKey_fu_138_statemt_we1),
    .statemt_d1(grp_AddRoundKey_fu_138_statemt_d1),
    .statemt_q1(statemt_q1),
    .n(grp_AddRoundKey_fu_138_n),
    .working_key(working_key)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_AddRoundKey_fu_138_ap_start_reg <= 1'b0;
    end else begin
      if((1'b1 == ap_CS_fsm_state10) | (exitcond6_fu_148_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
        grp_AddRoundKey_fu_138_ap_start_reg <= 1'b1;
      end else if(grp_AddRoundKey_fu_138_ap_ready == 1'b1) begin
        grp_AddRoundKey_fu_138_ap_start_reg <= 1'b0;
      end 
    end
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_ByteSub_ShiftRow_fu_131_ap_start_reg <= 1'b0;
    end else begin
      if((exitcond7_fu_165_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state5) | (exitcond7_fu_165_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state5)) begin
        grp_ByteSub_ShiftRow_fu_131_ap_start_reg <= 1'b1;
      end else if(grp_ByteSub_ShiftRow_fu_131_ap_ready == 1'b1) begin
        grp_ByteSub_ShiftRow_fu_131_ap_start_reg <= 1'b0;
      end 
    end
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_MixColumn_AddRoundKe_fu_122_ap_start_reg <= 1'b0;
    end else begin
      if(1'b1 == ap_CS_fsm_state7) begin
        grp_MixColumn_AddRoundKe_fu_122_ap_start_reg <= 1'b1;
      end else if(grp_MixColumn_AddRoundKe_fu_122_ap_ready == 1'b1) begin
        grp_MixColumn_AddRoundKe_fu_122_ap_start_reg <= 1'b0;
      end 
    end
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state4) & (grp_AddRoundKey_fu_138_ap_done == 1'b1)) begin
      if(working_key[2] == 1'b1) begin
        i_1_reg_99 <= temp100;
      end else begin
        i_1_reg_99 <= 4'd1;
      end
    end else if((grp_MixColumn_AddRoundKe_fu_122_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state8)) begin
      i_1_reg_99 <= i_4_reg_215;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state11) & (grp_AddRoundKey_fu_138_ap_done == 1'b1)) begin
      if(working_key[5] == 1'b1) begin
        i_2_reg_111 <= 6'd0;
      end else begin
        i_2_reg_111 <= temp104;
      end
    end else if(1'b1 == ap_CS_fsm_state13) begin
      i_2_reg_111 <= i_5_reg_223;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      i_reg_88 <= i_3_reg_197;
    end else if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      i_reg_88 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      i_3_reg_197 <= i_3_fu_154_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      i_4_reg_215 <= i_4_fu_171_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      i_5_reg_223 <= i_5_fu_183_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond_fu_177_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state12)) begin
      tmp_3_reg_228[5:0] <= tmp_3_fu_189_p1[5:0];
    end 
  end


  always @(posedge ap_clk) begin
    if((exitcond6_fu_148_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      tmp_reg_202[5:0] <= tmp_fu_160_p1[5:0];
    end 
  end


  always @(*) begin
    if((exitcond_fu_177_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state12)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if((exitcond_fu_177_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state12)) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      grp_AddRoundKey_fu_138_n = 6'd10;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      grp_AddRoundKey_fu_138_n = 6'd0;
    end else begin
      grp_AddRoundKey_fu_138_n = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      statemt1_address0 = tmp_3_reg_228;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt1_address0 = tmp_fu_160_p1;
    end else begin
      statemt1_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state13)) begin
      statemt1_ce0 = 1'b1;
    end else begin
      statemt1_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      statemt1_we0 = 1'b1;
    end else begin
      statemt1_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      statemt_address0 = tmp_3_fu_189_p1;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address0 = tmp_reg_202;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_address0 = grp_AddRoundKey_fu_138_statemt_address0;
    end else if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_address0 = grp_ByteSub_ShiftRow_fu_131_statemt_address0;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address0 = grp_MixColumn_AddRoundKe_fu_122_statemt_address0;
    end else begin
      statemt_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_address1 = grp_AddRoundKey_fu_138_statemt_address1;
    end else if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_address1 = grp_ByteSub_ShiftRow_fu_131_statemt_address1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address1 = grp_MixColumn_AddRoundKe_fu_122_statemt_address1;
    end else begin
      statemt_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state3)) begin
      statemt_ce0 = 1'b1;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_ce0 = grp_AddRoundKey_fu_138_statemt_ce0;
    end else if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_ce0 = grp_ByteSub_ShiftRow_fu_131_statemt_ce0;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_ce0 = grp_MixColumn_AddRoundKe_fu_122_statemt_ce0;
    end else begin
      statemt_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_ce1 = grp_AddRoundKey_fu_138_statemt_ce1;
    end else if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_ce1 = grp_ByteSub_ShiftRow_fu_131_statemt_ce1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_ce1 = grp_MixColumn_AddRoundKe_fu_122_statemt_ce1;
    end else begin
      statemt_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      statemt_d0 = statemt1_q0;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_d0 = grp_AddRoundKey_fu_138_statemt_d0;
    end else if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_d0 = grp_ByteSub_ShiftRow_fu_131_statemt_d0;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_d0 = grp_MixColumn_AddRoundKe_fu_122_statemt_d0;
    end else begin
      statemt_d0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_d1 = grp_AddRoundKey_fu_138_statemt_d1;
    end else if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_d1 = grp_ByteSub_ShiftRow_fu_131_statemt_d1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_d1 = grp_MixColumn_AddRoundKe_fu_122_statemt_d1;
    end else begin
      statemt_d1 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      statemt_we0 = 1'b1;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_we0 = grp_AddRoundKey_fu_138_statemt_we0;
    end else if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_we0 = grp_ByteSub_ShiftRow_fu_131_statemt_we0;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_we0 = grp_MixColumn_AddRoundKe_fu_122_statemt_we0;
    end else begin
      statemt_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_we1 = grp_AddRoundKey_fu_138_statemt_we1;
    end else if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_we1 = grp_ByteSub_ShiftRow_fu_131_statemt_we1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_we1 = grp_MixColumn_AddRoundKe_fu_122_statemt_we1;
    end else begin
      statemt_we1 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if((exitcond6_fu_148_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end
      end
      ap_ST_fsm_state3: begin
        ap_NS_fsm = ap_ST_fsm_state2;
      end
      ap_ST_fsm_state4: begin
        if((1'b1 == ap_CS_fsm_state4) & (grp_AddRoundKey_fu_138_ap_done == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end
      end
      ap_ST_fsm_state5: begin
        if((exitcond7_fu_165_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state5)) begin
          ap_NS_fsm = ap_ST_fsm_state9;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end
      end
      ap_ST_fsm_state6: begin
        if((1'b1 == ap_CS_fsm_state6) & (grp_ByteSub_ShiftRow_fu_131_ap_done == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end
      end
      ap_ST_fsm_state7: begin
        ap_NS_fsm = ap_ST_fsm_state8;
      end
      ap_ST_fsm_state8: begin
        if((grp_MixColumn_AddRoundKe_fu_122_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state8)) begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state9: begin
        if((1'b1 == ap_CS_fsm_state9) & (grp_ByteSub_ShiftRow_fu_131_ap_done == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state10;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state9;
        end
      end
      ap_ST_fsm_state10: begin
        ap_NS_fsm = ap_ST_fsm_state11;
      end
      ap_ST_fsm_state11: begin
        if((1'b1 == ap_CS_fsm_state11) & (grp_AddRoundKey_fu_138_ap_done == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state12;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state11;
        end
      end
      ap_ST_fsm_state12: begin
        if((exitcond_fu_177_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state12)) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state13;
        end
      end
      ap_ST_fsm_state13: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign exitcond6_fu_148_p2 = (i_reg_88 == 6'd32)? 1'b1 : 1'b0;
  assign exitcond7_fu_165_p2 = (i_1_reg_99 == 4'd10)? 1'b1 : 1'b0;
  assign exitcond_fu_177_p2 = (i_2_reg_111 == 6'd32)? 1'b1 : 1'b0;
  assign grp_AddRoundKey_fu_138_ap_start = grp_AddRoundKey_fu_138_ap_start_reg;
  assign grp_ByteSub_ShiftRow_fu_131_ap_start = grp_ByteSub_ShiftRow_fu_131_ap_start_reg;
  assign grp_MixColumn_AddRoundKe_fu_122_ap_start = grp_MixColumn_AddRoundKe_fu_122_ap_start_reg;
  assign i_3_fu_154_p2 = i_reg_88 + 6'd1;
  assign i_4_fu_171_p2 = i_1_reg_99 + 4'd1;
  assign i_5_fu_183_p2 = i_2_reg_111 + 6'd1;
  assign statemt1_d0 = statemt_q0;
  assign tmp_3_fu_189_p1 = i_2_reg_111;
  assign tmp_fu_160_p1 = i_reg_88;

  always @(posedge ap_clk) begin
    tmp_reg_202[63:6] <= 58'b0000000000000000000000000000000000000000000000000000000000;
    tmp_3_reg_228[63:6] <= 58'b0000000000000000000000000000000000000000000000000000000000;
  end

  assign temp100 = temp102 * temp103;
  assign temp103 = (working_key[0] == 1'b1)? grp_AddRoundKey_fu_138_statemt_ce0 + ap_CS_fsm_state2 : grp_MixColumn_AddRoundKe_fu_122_statemt_d0 + grp_ByteSub_ShiftRow_fu_131_ap_idle;
  assign temp102 = (working_key[1] == 1'b1)? grp_ByteSub_ShiftRow_fu_131_ap_done + grp_AddRoundKey_fu_138_ap_done : ap_CS_fsm_state1 + statemt_q1;
  assign temp104 = temp106 * temp107;
  assign temp107 = (working_key[3] == 1'b1)? grp_ByteSub_ShiftRow_fu_131_statemt_we1 + ap_CS_fsm_state13 : grp_MixColumn_AddRoundKe_fu_122_statemt_we1 + grp_AddRoundKey_fu_138_statemt_d1;
  assign temp106 = (working_key[4] == 1'b1)? grp_ByteSub_ShiftRow_fu_131_statemt_address1 + grp_ByteSub_ShiftRow_fu_131_statemt_d1 : grp_AddRoundKey_fu_138_statemt_we1 + ap_CS_fsm_state11;

endmodule



module decode
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  input_r,
  ih_i,
  ih_o,
  ih_o_ap_vld,
  dec_del_bpl_address0,
  dec_del_bpl_ce0,
  dec_del_bpl_we0,
  dec_del_bpl_d0,
  dec_del_bpl_q0,
  dec_del_dltx_address0,
  dec_del_dltx_ce0,
  dec_del_dltx_we0,
  dec_del_dltx_d0,
  dec_del_dltx_q0,
  dec_del_dltx_address1,
  dec_del_dltx_ce1,
  dec_del_dltx_we1,
  dec_del_dltx_d1,
  dec_del_dltx_q1,
  dec_rlt1_i,
  dec_rlt1_o,
  dec_rlt1_o_ap_vld,
  dec_al1_i,
  dec_al1_o,
  dec_al1_o_ap_vld,
  dec_rlt2_i,
  dec_rlt2_o,
  dec_rlt2_o_ap_vld,
  dec_al2_i,
  dec_al2_o,
  dec_al2_o_ap_vld,
  dec_detl_i,
  dec_detl_o,
  dec_detl_o_ap_vld,
  il,
  dec_nbl_i,
  dec_nbl_o,
  dec_nbl_o_ap_vld,
  dec_plt1_i,
  dec_plt1_o,
  dec_plt1_o_ap_vld,
  dec_plt2_i,
  dec_plt2_o,
  dec_plt2_o_ap_vld,
  dec_del_bph_address0,
  dec_del_bph_ce0,
  dec_del_bph_we0,
  dec_del_bph_d0,
  dec_del_bph_q0,
  dec_del_dhx_address0,
  dec_del_dhx_ce0,
  dec_del_dhx_we0,
  dec_del_dhx_d0,
  dec_del_dhx_q0,
  dec_del_dhx_address1,
  dec_del_dhx_ce1,
  dec_del_dhx_we1,
  dec_del_dhx_d1,
  dec_del_dhx_q1,
  dec_rh1_i,
  dec_rh1_o,
  dec_rh1_o_ap_vld,
  dec_ah1_i,
  dec_ah1_o,
  dec_ah1_o_ap_vld,
  dec_rh2_i,
  dec_rh2_o,
  dec_rh2_o_ap_vld,
  dec_ah2_i,
  dec_ah2_o,
  dec_ah2_o_ap_vld,
  dec_deth_i,
  dec_deth_o,
  dec_deth_o_ap_vld,
  dec_nbh_i,
  dec_nbh_o,
  dec_nbh_o_ap_vld,
  dec_ph1_i,
  dec_ph1_o,
  dec_ph1_o_ap_vld,
  dec_ph2_i,
  dec_ph2_o,
  dec_ph2_o_ap_vld,
  accumc_address0,
  accumc_ce0,
  accumc_we0,
  accumc_d0,
  accumc_q0,
  accumd_address0,
  accumd_ce0,
  accumd_we0,
  accumd_d0,
  accumd_q0
);

  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  input [31:0] input_r;
  input [31:0] ih_i;
  output [31:0] ih_o;
  output ih_o_ap_vld;
  output [2:0] dec_del_bpl_address0;
  output dec_del_bpl_ce0;
  output dec_del_bpl_we0;
  output [31:0] dec_del_bpl_d0;
  input [31:0] dec_del_bpl_q0;
  output [2:0] dec_del_dltx_address0;
  output dec_del_dltx_ce0;
  output dec_del_dltx_we0;
  output [31:0] dec_del_dltx_d0;
  input [31:0] dec_del_dltx_q0;
  output [2:0] dec_del_dltx_address1;
  output dec_del_dltx_ce1;
  output dec_del_dltx_we1;
  output [31:0] dec_del_dltx_d1;
  input [31:0] dec_del_dltx_q1;
  input [31:0] dec_rlt1_i;
  output [31:0] dec_rlt1_o;
  output dec_rlt1_o_ap_vld;
  input [31:0] dec_al1_i;
  output [31:0] dec_al1_o;
  output dec_al1_o_ap_vld;
  input [31:0] dec_rlt2_i;
  output [31:0] dec_rlt2_o;
  output dec_rlt2_o_ap_vld;
  input [31:0] dec_al2_i;
  output [31:0] dec_al2_o;
  output dec_al2_o_ap_vld;
  input [14:0] dec_detl_i;
  output [14:0] dec_detl_o;
  output dec_detl_o_ap_vld;
  input [5:0] il;
  input [31:0] dec_nbl_i;
  output [31:0] dec_nbl_o;
  output dec_nbl_o_ap_vld;
  input [31:0] dec_plt1_i;
  output [31:0] dec_plt1_o;
  output dec_plt1_o_ap_vld;
  input [31:0] dec_plt2_i;
  output [31:0] dec_plt2_o;
  output dec_plt2_o_ap_vld;
  output [2:0] dec_del_bph_address0;
  output dec_del_bph_ce0;
  output dec_del_bph_we0;
  output [31:0] dec_del_bph_d0;
  input [31:0] dec_del_bph_q0;
  output [2:0] dec_del_dhx_address0;
  output dec_del_dhx_ce0;
  output dec_del_dhx_we0;
  output [31:0] dec_del_dhx_d0;
  input [31:0] dec_del_dhx_q0;
  output [2:0] dec_del_dhx_address1;
  output dec_del_dhx_ce1;
  output dec_del_dhx_we1;
  output [31:0] dec_del_dhx_d1;
  input [31:0] dec_del_dhx_q1;
  input [31:0] dec_rh1_i;
  output [31:0] dec_rh1_o;
  output dec_rh1_o_ap_vld;
  input [31:0] dec_ah1_i;
  output [31:0] dec_ah1_o;
  output dec_ah1_o_ap_vld;
  input [31:0] dec_rh2_i;
  output [31:0] dec_rh2_o;
  output dec_rh2_o_ap_vld;
  input [31:0] dec_ah2_i;
  output [31:0] dec_ah2_o;
  output dec_ah2_o_ap_vld;
  input [14:0] dec_deth_i;
  output [14:0] dec_deth_o;
  output dec_deth_o_ap_vld;
  input [31:0] dec_nbh_i;
  output [31:0] dec_nbh_o;
  output dec_nbh_o_ap_vld;
  input [31:0] dec_ph1_i;
  output [31:0] dec_ph1_o;
  output dec_ph1_o_ap_vld;
  input [31:0] dec_ph2_i;
  output [31:0] dec_ph2_o;
  output dec_ph2_o_ap_vld;
  output [3:0] accumc_address0;
  output accumc_ce0;
  output accumc_we0;
  output [31:0] accumc_d0;
  input [31:0] accumc_q0;
  output [3:0] accumd_address0;
  output accumd_ce0;
  output accumd_we0;
  output [31:0] accumd_d0;
  input [31:0] accumd_q0;

  decode_0_obf
  i0
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .input_r(input_r),
    .ih_i(ih_i),
    .ih_o(ih_o),
    .ih_o_ap_vld(ih_o_ap_vld),
    .dec_del_bpl_address0(dec_del_bpl_address0),
    .dec_del_bpl_ce0(dec_del_bpl_ce0),
    .dec_del_bpl_we0(dec_del_bpl_we0),
    .dec_del_bpl_d0(dec_del_bpl_d0),
    .dec_del_bpl_q0(dec_del_bpl_q0),
    .dec_del_dltx_address0(dec_del_dltx_address0),
    .dec_del_dltx_ce0(dec_del_dltx_ce0),
    .dec_del_dltx_we0(dec_del_dltx_we0),
    .dec_del_dltx_d0(dec_del_dltx_d0),
    .dec_del_dltx_q0(dec_del_dltx_q0),
    .dec_del_dltx_address1(dec_del_dltx_address1),
    .dec_del_dltx_ce1(dec_del_dltx_ce1),
    .dec_del_dltx_we1(dec_del_dltx_we1),
    .dec_del_dltx_d1(dec_del_dltx_d1),
    .dec_del_dltx_q1(dec_del_dltx_q1),
    .dec_rlt1_i(dec_rlt1_i),
    .dec_rlt1_o(dec_rlt1_o),
    .dec_rlt1_o_ap_vld(dec_rlt1_o_ap_vld),
    .dec_al1_i(dec_al1_i),
    .dec_al1_o(dec_al1_o),
    .dec_al1_o_ap_vld(dec_al1_o_ap_vld),
    .dec_rlt2_i(dec_rlt2_i),
    .dec_rlt2_o(dec_rlt2_o),
    .dec_rlt2_o_ap_vld(dec_rlt2_o_ap_vld),
    .dec_al2_i(dec_al2_i),
    .dec_al2_o(dec_al2_o),
    .dec_al2_o_ap_vld(dec_al2_o_ap_vld),
    .dec_detl_i(dec_detl_i),
    .dec_detl_o(dec_detl_o),
    .dec_detl_o_ap_vld(dec_detl_o_ap_vld),
    .il(il),
    .dec_nbl_i(dec_nbl_i),
    .dec_nbl_o(dec_nbl_o),
    .dec_nbl_o_ap_vld(dec_nbl_o_ap_vld),
    .dec_plt1_i(dec_plt1_i),
    .dec_plt1_o(dec_plt1_o),
    .dec_plt1_o_ap_vld(dec_plt1_o_ap_vld),
    .dec_plt2_i(dec_plt2_i),
    .dec_plt2_o(dec_plt2_o),
    .dec_plt2_o_ap_vld(dec_plt2_o_ap_vld),
    .dec_del_bph_address0(dec_del_bph_address0),
    .dec_del_bph_ce0(dec_del_bph_ce0),
    .dec_del_bph_we0(dec_del_bph_we0),
    .dec_del_bph_d0(dec_del_bph_d0),
    .dec_del_bph_q0(dec_del_bph_q0),
    .dec_del_dhx_address0(dec_del_dhx_address0),
    .dec_del_dhx_ce0(dec_del_dhx_ce0),
    .dec_del_dhx_we0(dec_del_dhx_we0),
    .dec_del_dhx_d0(dec_del_dhx_d0),
    .dec_del_dhx_q0(dec_del_dhx_q0),
    .dec_del_dhx_address1(dec_del_dhx_address1),
    .dec_del_dhx_ce1(dec_del_dhx_ce1),
    .dec_del_dhx_we1(dec_del_dhx_we1),
    .dec_del_dhx_d1(dec_del_dhx_d1),
    .dec_del_dhx_q1(dec_del_dhx_q1),
    .dec_rh1_i(dec_rh1_i),
    .dec_rh1_o(dec_rh1_o),
    .dec_rh1_o_ap_vld(dec_rh1_o_ap_vld),
    .dec_ah1_i(dec_ah1_i),
    .dec_ah1_o(dec_ah1_o),
    .dec_ah1_o_ap_vld(dec_ah1_o_ap_vld),
    .dec_rh2_i(dec_rh2_i),
    .dec_rh2_o(dec_rh2_o),
    .dec_rh2_o_ap_vld(dec_rh2_o_ap_vld),
    .dec_ah2_i(dec_ah2_i),
    .dec_ah2_o(dec_ah2_o),
    .dec_ah2_o_ap_vld(dec_ah2_o_ap_vld),
    .dec_deth_i(dec_deth_i),
    .dec_deth_o(dec_deth_o),
    .dec_deth_o_ap_vld(dec_deth_o_ap_vld),
    .dec_nbh_i(dec_nbh_i),
    .dec_nbh_o(dec_nbh_o),
    .dec_nbh_o_ap_vld(dec_nbh_o_ap_vld),
    .dec_ph1_i(dec_ph1_i),
    .dec_ph1_o(dec_ph1_o),
    .dec_ph1_o_ap_vld(dec_ph1_o_ap_vld),
    .dec_ph2_i(dec_ph2_i),
    .dec_ph2_o(dec_ph2_o),
    .dec_ph2_o_ap_vld(dec_ph2_o_ap_vld),
    .accumc_address0(accumc_address0),
    .accumc_ce0(accumc_ce0),
    .accumc_we0(accumc_we0),
    .accumc_d0(accumc_d0),
    .accumc_q0(accumc_q0),
    .accumd_address0(accumd_address0),
    .accumd_ce0(accumd_ce0),
    .accumd_we0(accumd_we0),
    .accumd_d0(accumd_d0),
    .accumd_q0(accumd_q0),
    .working_key(12287'b11001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101010100110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101010100110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101010100110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101010100110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101010100110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101010100110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101010100110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101010100110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101111111101100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010011001010101010101010101010000010101010101010101010010101011111110100110101010010010101101010101110100110101010010010101101011110110010101010101010101010100000101010101010101010100101010111111101001101010100100101011010101011101001101010100100101011010101001100101010101010101010101000001010101010101010101001010101111111010011010101001001010110101010111010011010101001001010110101010)
  );


endmodule


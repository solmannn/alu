
module backprop_0_obf
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  weights_address0,
  weights_ce0,
  weights_we0,
  weights_d0,
  weights_q0,
  inputs_address0,
  inputs_ce0,
  inputs_q0,
  targets_address0,
  targets_ce0,
  targets_q0,
  locking_key
);

  parameter ap_ST_fsm_state1 = 201'd1;
  parameter ap_ST_fsm_state2 = 201'd2;
  parameter ap_ST_fsm_state3 = 201'd4;
  parameter ap_ST_fsm_state4 = 201'd8;
  parameter ap_ST_fsm_state5 = 201'd16;
  parameter ap_ST_fsm_state6 = 201'd32;
  parameter ap_ST_fsm_state7 = 201'd64;
  parameter ap_ST_fsm_state8 = 201'd128;
  parameter ap_ST_fsm_state9 = 201'd256;
  parameter ap_ST_fsm_state10 = 201'd512;
  parameter ap_ST_fsm_state11 = 201'd1024;
  parameter ap_ST_fsm_state12 = 201'd2048;
  parameter ap_ST_fsm_state13 = 201'd4096;
  parameter ap_ST_fsm_state14 = 201'd8192;
  parameter ap_ST_fsm_state15 = 201'd16384;
  parameter ap_ST_fsm_state16 = 201'd32768;
  parameter ap_ST_fsm_state17 = 201'd65536;
  parameter ap_ST_fsm_state18 = 201'd131072;
  parameter ap_ST_fsm_state19 = 201'd262144;
  parameter ap_ST_fsm_state20 = 201'd524288;
  parameter ap_ST_fsm_state21 = 201'd1048576;
  parameter ap_ST_fsm_state22 = 201'd2097152;
  parameter ap_ST_fsm_state23 = 201'd4194304;
  parameter ap_ST_fsm_state24 = 201'd8388608;
  parameter ap_ST_fsm_state25 = 201'd16777216;
  parameter ap_ST_fsm_state26 = 201'd33554432;
  parameter ap_ST_fsm_state27 = 201'd67108864;
  parameter ap_ST_fsm_state28 = 201'd134217728;
  parameter ap_ST_fsm_state29 = 201'd268435456;
  parameter ap_ST_fsm_state30 = 201'd536870912;
  parameter ap_ST_fsm_state31 = 201'd1073741824;
  parameter ap_ST_fsm_state32 = 201'd2147483648;
  parameter ap_ST_fsm_state33 = 201'd4294967296;
  parameter ap_ST_fsm_state34 = 201'd8589934592;
  parameter ap_ST_fsm_state35 = 201'd17179869184;
  parameter ap_ST_fsm_state36 = 201'd34359738368;
  parameter ap_ST_fsm_state37 = 201'd68719476736;
  parameter ap_ST_fsm_state38 = 201'd137438953472;
  parameter ap_ST_fsm_state39 = 201'd274877906944;
  parameter ap_ST_fsm_state40 = 201'd549755813888;
  parameter ap_ST_fsm_state41 = 201'd1099511627776;
  parameter ap_ST_fsm_state42 = 201'd2199023255552;
  parameter ap_ST_fsm_state43 = 201'd4398046511104;
  parameter ap_ST_fsm_state44 = 201'd8796093022208;
  parameter ap_ST_fsm_state45 = 201'd17592186044416;
  parameter ap_ST_fsm_state46 = 201'd35184372088832;
  parameter ap_ST_fsm_state47 = 201'd70368744177664;
  parameter ap_ST_fsm_state48 = 201'd140737488355328;
  parameter ap_ST_fsm_state49 = 201'd281474976710656;
  parameter ap_ST_fsm_state50 = 201'd562949953421312;
  parameter ap_ST_fsm_state51 = 201'd1125899906842624;
  parameter ap_ST_fsm_state52 = 201'd2251799813685248;
  parameter ap_ST_fsm_state53 = 201'd4503599627370496;
  parameter ap_ST_fsm_state54 = 201'd9007199254740992;
  parameter ap_ST_fsm_state55 = 201'd18014398509481984;
  parameter ap_ST_fsm_state56 = 201'd36028797018963968;
  parameter ap_ST_fsm_state57 = 201'd72057594037927936;
  parameter ap_ST_fsm_state58 = 201'd144115188075855872;
  parameter ap_ST_fsm_state59 = 201'd288230376151711744;
  parameter ap_ST_fsm_state60 = 201'd576460752303423488;
  parameter ap_ST_fsm_state61 = 201'd1152921504606846976;
  parameter ap_ST_fsm_state62 = 201'd2305843009213693952;
  parameter ap_ST_fsm_state63 = 201'd4611686018427387904;
  parameter ap_ST_fsm_state64 = 201'd9223372036854775808;
  parameter ap_ST_fsm_state65 = 201'd18446744073709551616;
  parameter ap_ST_fsm_state66 = 201'd36893488147419103232;
  parameter ap_ST_fsm_state67 = 201'd73786976294838206464;
  parameter ap_ST_fsm_state68 = 201'd147573952589676412928;
  parameter ap_ST_fsm_state69 = 201'd295147905179352825856;
  parameter ap_ST_fsm_state70 = 201'd590295810358705651712;
  parameter ap_ST_fsm_state71 = 201'd1180591620717411303424;
  parameter ap_ST_fsm_state72 = 201'd2361183241434822606848;
  parameter ap_ST_fsm_state73 = 201'd4722366482869645213696;
  parameter ap_ST_fsm_state74 = 201'd9444732965739290427392;
  parameter ap_ST_fsm_state75 = 201'd18889465931478580854784;
  parameter ap_ST_fsm_state76 = 201'd37778931862957161709568;
  parameter ap_ST_fsm_state77 = 201'd75557863725914323419136;
  parameter ap_ST_fsm_state78 = 201'd151115727451828646838272;
  parameter ap_ST_fsm_state79 = 201'd302231454903657293676544;
  parameter ap_ST_fsm_state80 = 201'd604462909807314587353088;
  parameter ap_ST_fsm_state81 = 201'd1208925819614629174706176;
  parameter ap_ST_fsm_state82 = 201'd2417851639229258349412352;
  parameter ap_ST_fsm_state83 = 201'd4835703278458516698824704;
  parameter ap_ST_fsm_state84 = 201'd9671406556917033397649408;
  parameter ap_ST_fsm_state85 = 201'd19342813113834066795298816;
  parameter ap_ST_fsm_state86 = 201'd38685626227668133590597632;
  parameter ap_ST_fsm_state87 = 201'd77371252455336267181195264;
  parameter ap_ST_fsm_state88 = 201'd154742504910672534362390528;
  parameter ap_ST_fsm_state89 = 201'd309485009821345068724781056;
  parameter ap_ST_fsm_state90 = 201'd618970019642690137449562112;
  parameter ap_ST_fsm_state91 = 201'd1237940039285380274899124224;
  parameter ap_ST_fsm_state92 = 201'd2475880078570760549798248448;
  parameter ap_ST_fsm_state93 = 201'd4951760157141521099596496896;
  parameter ap_ST_fsm_state94 = 201'd9903520314283042199192993792;
  parameter ap_ST_fsm_state95 = 201'd19807040628566084398385987584;
  parameter ap_ST_fsm_state96 = 201'd39614081257132168796771975168;
  parameter ap_ST_fsm_state97 = 201'd79228162514264337593543950336;
  parameter ap_ST_fsm_state98 = 201'd158456325028528675187087900672;
  parameter ap_ST_fsm_state99 = 201'd316912650057057350374175801344;
  parameter ap_ST_fsm_state100 = 201'd633825300114114700748351602688;
  parameter ap_ST_fsm_state101 = 201'd1267650600228229401496703205376;
  parameter ap_ST_fsm_state102 = 201'd2535301200456458802993406410752;
  parameter ap_ST_fsm_state103 = 201'd5070602400912917605986812821504;
  parameter ap_ST_fsm_state104 = 201'd10141204801825835211973625643008;
  parameter ap_ST_fsm_state105 = 201'd20282409603651670423947251286016;
  parameter ap_ST_fsm_state106 = 201'd40564819207303340847894502572032;
  parameter ap_ST_fsm_state107 = 201'd81129638414606681695789005144064;
  parameter ap_ST_fsm_state108 = 201'd162259276829213363391578010288128;
  parameter ap_ST_fsm_state109 = 201'd324518553658426726783156020576256;
  parameter ap_ST_fsm_state110 = 201'd649037107316853453566312041152512;
  parameter ap_ST_fsm_state111 = 201'd1298074214633706907132624082305024;
  parameter ap_ST_fsm_state112 = 201'd2596148429267413814265248164610048;
  parameter ap_ST_fsm_state113 = 201'd5192296858534827628530496329220096;
  parameter ap_ST_fsm_state114 = 201'd10384593717069655257060992658440192;
  parameter ap_ST_fsm_state115 = 201'd20769187434139310514121985316880384;
  parameter ap_ST_fsm_state116 = 201'd41538374868278621028243970633760768;
  parameter ap_ST_fsm_state117 = 201'd83076749736557242056487941267521536;
  parameter ap_ST_fsm_state118 = 201'd166153499473114484112975882535043072;
  parameter ap_ST_fsm_state119 = 201'd332306998946228968225951765070086144;
  parameter ap_ST_fsm_state120 = 201'd664613997892457936451903530140172288;
  parameter ap_ST_fsm_state121 = 201'd1329227995784915872903807060280344576;
  parameter ap_ST_fsm_state122 = 201'd2658455991569831745807614120560689152;
  parameter ap_ST_fsm_state123 = 201'd5316911983139663491615228241121378304;
  parameter ap_ST_fsm_state124 = 201'd10633823966279326983230456482242756608;
  parameter ap_ST_fsm_state125 = 201'd21267647932558653966460912964485513216;
  parameter ap_ST_fsm_state126 = 201'd42535295865117307932921825928971026432;
  parameter ap_ST_fsm_state127 = 201'd85070591730234615865843651857942052864;
  parameter ap_ST_fsm_state128 = 201'd170141183460469231731687303715884105728;
  parameter ap_ST_fsm_state129 = 201'd340282366920938463463374607431768211456;
  parameter ap_ST_fsm_state130 = 201'd680564733841876926926749214863536422912;
  parameter ap_ST_fsm_state131 = 201'd1361129467683753853853498429727072845824;
  parameter ap_ST_fsm_state132 = 201'd2722258935367507707706996859454145691648;
  parameter ap_ST_fsm_state133 = 201'd5444517870735015415413993718908291383296;
  parameter ap_ST_fsm_state134 = 201'd10889035741470030830827987437816582766592;
  parameter ap_ST_fsm_state135 = 201'd21778071482940061661655974875633165533184;
  parameter ap_ST_fsm_state136 = 201'd43556142965880123323311949751266331066368;
  parameter ap_ST_fsm_state137 = 201'd87112285931760246646623899502532662132736;
  parameter ap_ST_fsm_state138 = 201'd174224571863520493293247799005065324265472;
  parameter ap_ST_fsm_state139 = 201'd348449143727040986586495598010130648530944;
  parameter ap_ST_fsm_state140 = 201'd696898287454081973172991196020261297061888;
  parameter ap_ST_fsm_state141 = 201'd1393796574908163946345982392040522594123776;
  parameter ap_ST_fsm_state142 = 201'd2787593149816327892691964784081045188247552;
  parameter ap_ST_fsm_state143 = 201'd5575186299632655785383929568162090376495104;
  parameter ap_ST_fsm_state144 = 201'd11150372599265311570767859136324180752990208;
  parameter ap_ST_fsm_state145 = 201'd22300745198530623141535718272648361505980416;
  parameter ap_ST_fsm_state146 = 201'd44601490397061246283071436545296723011960832;
  parameter ap_ST_fsm_state147 = 201'd89202980794122492566142873090593446023921664;
  parameter ap_ST_fsm_state148 = 201'd178405961588244985132285746181186892047843328;
  parameter ap_ST_fsm_state149 = 201'd356811923176489970264571492362373784095686656;
  parameter ap_ST_fsm_state150 = 201'd713623846352979940529142984724747568191373312;
  parameter ap_ST_fsm_state151 = 201'd1427247692705959881058285969449495136382746624;
  parameter ap_ST_fsm_state152 = 201'd2854495385411919762116571938898990272765493248;
  parameter ap_ST_fsm_state153 = 201'd5708990770823839524233143877797980545530986496;
  parameter ap_ST_fsm_state154 = 201'd11417981541647679048466287755595961091061972992;
  parameter ap_ST_fsm_state155 = 201'd22835963083295358096932575511191922182123945984;
  parameter ap_ST_fsm_state156 = 201'd45671926166590716193865151022383844364247891968;
  parameter ap_ST_fsm_state157 = 201'd91343852333181432387730302044767688728495783936;
  parameter ap_ST_fsm_state158 = 201'd182687704666362864775460604089535377456991567872;
  parameter ap_ST_fsm_state159 = 201'd365375409332725729550921208179070754913983135744;
  parameter ap_ST_fsm_state160 = 201'd730750818665451459101842416358141509827966271488;
  parameter ap_ST_fsm_state161 = 201'd1461501637330902918203684832716283019655932542976;
  parameter ap_ST_fsm_state162 = 201'd2923003274661805836407369665432566039311865085952;
  parameter ap_ST_fsm_state163 = 201'd5846006549323611672814739330865132078623730171904;
  parameter ap_ST_fsm_state164 = 201'd11692013098647223345629478661730264157247460343808;
  parameter ap_ST_fsm_state165 = 201'd23384026197294446691258957323460528314494920687616;
  parameter ap_ST_fsm_state166 = 201'd46768052394588893382517914646921056628989841375232;
  parameter ap_ST_fsm_state167 = 201'd93536104789177786765035829293842113257979682750464;
  parameter ap_ST_fsm_state168 = 201'd187072209578355573530071658587684226515959365500928;
  parameter ap_ST_fsm_state169 = 201'd374144419156711147060143317175368453031918731001856;
  parameter ap_ST_fsm_state170 = 201'd748288838313422294120286634350736906063837462003712;
  parameter ap_ST_fsm_state171 = 201'd1496577676626844588240573268701473812127674924007424;
  parameter ap_ST_fsm_state172 = 201'd2993155353253689176481146537402947624255349848014848;
  parameter ap_ST_fsm_state173 = 201'd5986310706507378352962293074805895248510699696029696;
  parameter ap_ST_fsm_state174 = 201'd11972621413014756705924586149611790497021399392059392;
  parameter ap_ST_fsm_state175 = 201'd23945242826029513411849172299223580994042798784118784;
  parameter ap_ST_fsm_state176 = 201'd47890485652059026823698344598447161988085597568237568;
  parameter ap_ST_fsm_state177 = 201'd95780971304118053647396689196894323976171195136475136;
  parameter ap_ST_fsm_state178 = 201'd191561942608236107294793378393788647952342390272950272;
  parameter ap_ST_fsm_state179 = 201'd383123885216472214589586756787577295904684780545900544;
  parameter ap_ST_fsm_state180 = 201'd766247770432944429179173513575154591809369561091801088;
  parameter ap_ST_fsm_state181 = 201'd1532495540865888858358347027150309183618739122183602176;
  parameter ap_ST_fsm_state182 = 201'd3064991081731777716716694054300618367237478244367204352;
  parameter ap_ST_fsm_state183 = 201'd6129982163463555433433388108601236734474956488734408704;
  parameter ap_ST_fsm_state184 = 201'd12259964326927110866866776217202473468949912977468817408;
  parameter ap_ST_fsm_state185 = 201'd24519928653854221733733552434404946937899825954937634816;
  parameter ap_ST_fsm_state186 = 201'd49039857307708443467467104868809893875799651909875269632;
  parameter ap_ST_fsm_state187 = 201'd98079714615416886934934209737619787751599303819750539264;
  parameter ap_ST_fsm_state188 = 201'd196159429230833773869868419475239575503198607639501078528;
  parameter ap_ST_fsm_state189 = 201'd392318858461667547739736838950479151006397215279002157056;
  parameter ap_ST_fsm_state190 = 201'd784637716923335095479473677900958302012794430558004314112;
  parameter ap_ST_fsm_state191 = 201'd1569275433846670190958947355801916604025588861116008628224;
  parameter ap_ST_fsm_state192 = 201'd3138550867693340381917894711603833208051177722232017256448;
  parameter ap_ST_fsm_state193 = 201'd6277101735386680763835789423207666416102355444464034512896;
  parameter ap_ST_fsm_state194 = 201'd12554203470773361527671578846415332832204710888928069025792;
  parameter ap_ST_fsm_state195 = 201'd25108406941546723055343157692830665664409421777856138051584;
  parameter ap_ST_fsm_state196 = 201'd50216813883093446110686315385661331328818843555712276103168;
  parameter ap_ST_fsm_state197 = 201'd100433627766186892221372630771322662657637687111424552206336;
  parameter ap_ST_fsm_state198 = 201'd200867255532373784442745261542645325315275374222849104412672;
  parameter ap_ST_fsm_state199 = 201'd401734511064747568885490523085290650630550748445698208825344;
  parameter ap_ST_fsm_state200 = 201'd803469022129495137770981046170581301261101496891396417650688;
  parameter ap_ST_fsm_state201 = 201'd1606938044258990275541962092341162602522202993782792835301376;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [7:0] weights_address0;
  output weights_ce0;
  output weights_we0;
  output [63:0] weights_d0;
  input [63:0] weights_q0;
  output [8:0] inputs_address0;
  output inputs_ce0;
  input [63:0] inputs_q0;
  output [9:0] targets_address0;
  output targets_ce0;
  input [63:0] targets_q0;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [7:0] weights_address0;
  reg weights_ce0;
  reg weights_we0;
  reg inputs_ce0;
  reg targets_ce0;
  reg [200:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  wire [63:0] activations_q0;
  reg [63:0] reg_583;
  wire ap_CS_fsm_state14;
  wire ap_CS_fsm_state69;
  wire ap_CS_fsm_state178;
  reg [63:0] reg_590;
  wire ap_CS_fsm_state118;
  wire ap_CS_fsm_state190;
  wire [63:0] grp_fu_566_p2;
  reg [63:0] reg_596;
  wire ap_CS_fsm_state19;
  wire ap_CS_fsm_state114;
  wire ap_CS_fsm_state123;
  wire ap_CS_fsm_state174;
  wire ap_CS_fsm_state185;
  wire ap_CS_fsm_state195;
  wire [63:0] grp_fu_578_p2;
  reg [63:0] reg_604;
  wire ap_CS_fsm_state37;
  wire ap_CS_fsm_state82;
  wire ap_CS_fsm_state142;
  wire [63:0] grp_fu_559_p2;
  reg [63:0] reg_609;
  wire ap_CS_fsm_state42;
  wire ap_CS_fsm_state74;
  wire ap_CS_fsm_state147;
  wire ap_CS_fsm_state200;
  wire [63:0] grp_fu_573_p2;
  reg [63:0] reg_617;
  wire ap_CS_fsm_state64;
  wire ap_CS_fsm_state109;
  wire ap_CS_fsm_state169;
  wire [63:0] deltas_q0;
  reg [63:0] reg_623;
  wire ap_CS_fsm_state180;
  wire [1:0] ee_fu_634_p2;
  reg [1:0] ee_reg_1581;
  wire ap_CS_fsm_state2;
  wire [5:0] add_ln160_fu_664_p2;
  reg [5:0] add_ln160_reg_1586;
  wire [0:0] icmp_ln156_fu_628_p2;
  wire [3:0] rows_fu_676_p2;
  reg [3:0] rows_reg_1594;
  wire ap_CS_fsm_state3;
  wire [9:0] add_ln160_2_fu_720_p2;
  reg [9:0] add_ln160_2_reg_1599;
  wire [0:0] icmp_ln157_fu_670_p2;
  wire [3:0] cols_fu_732_p2;
  wire ap_CS_fsm_state4;
  wire [6:0] ee_2_fu_758_p2;
  reg [6:0] ee_2_reg_1615;
  wire ap_CS_fsm_state5;
  wire [6:0] jj_1_fu_770_p2;
  reg [6:0] jj_1_reg_1623;
  wire ap_CS_fsm_state6;
  wire [1:0] cols_2_fu_782_p2;
  reg [1:0] cols_2_reg_1631;
  wire ap_CS_fsm_state7;
  wire [5:0] add_ln170_fu_812_p2;
  reg [5:0] add_ln170_reg_1636;
  wire [0:0] icmp_ln168_fu_776_p2;
  wire [9:0] zext_ln52_fu_826_p1;
  reg [9:0] zext_ln52_reg_1641;
  wire [10:0] add_ln52_fu_854_p2;
  reg [10:0] add_ln52_reg_1646;
  wire [3:0] rows_2_fu_866_p2;
  wire ap_CS_fsm_state8;
  wire [2:0] i_fu_892_p2;
  reg [2:0] i_reg_1662;
  wire ap_CS_fsm_state9;
  wire [0:0] icmp_ln34_fu_886_p2;
  wire [1:0] i_1_fu_923_p2;
  reg [1:0] i_1_reg_1675;
  wire ap_CS_fsm_state11;
  wire [5:0] add_ln21_fu_953_p2;
  reg [5:0] add_ln21_reg_1680;
  wire [0:0] icmp_ln39_fu_917_p2;
  wire [3:0] select_ln40_fu_963_p3;
  reg [3:0] select_ln40_reg_1685;
  wire [5:0] add_ln23_fu_995_p2;
  reg [5:0] add_ln23_reg_1690;
  wire [3:0] ii_fu_1007_p2;
  reg [3:0] ii_reg_1698;
  wire ap_CS_fsm_state12;
  wire [8:0] zext_ln23_2_fu_1013_p1;
  reg [8:0] zext_ln23_2_reg_1703;
  wire [0:0] icmp_ln18_fu_1001_p2;
  reg [4:0] activations_addr_5_reg_1708;
  wire [3:0] jj_fu_1036_p2;
  reg [3:0] jj_reg_1716;
  wire ap_CS_fsm_state13;
  wire [0:0] icmp_ln20_fu_1031_p2;
  wire [63:0] xor_ln7_1_fu_1096_p2;
  reg [63:0] xor_ln7_1_reg_1731;
  wire ap_CS_fsm_state24;
  wire [63:0] bitcast_ln7_3_fu_1102_p1;
  wire ap_CS_fsm_state25;
  wire [1:0] i_3_fu_1112_p2;
  reg [1:0] i_3_reg_1749;
  wire ap_CS_fsm_state66;
  wire [5:0] add_ln112_fu_1142_p2;
  reg [5:0] add_ln112_reg_1754;
  wire [0:0] icmp_ln110_fu_1106_p2;
  wire [3:0] j_fu_1154_p2;
  wire ap_CS_fsm_state67;
  wire [3:0] i_2_fu_1180_p2;
  reg [3:0] i_2_reg_1770;
  wire ap_CS_fsm_state68;
  wire [4:0] zext_ln52_3_fu_1186_p1;
  reg [4:0] zext_ln52_3_reg_1775;
  wire [0:0] icmp_ln51_fu_1174_p2;
  reg [63:0] targets_load_reg_1790;
  wire [63:0] xor_ln7_fu_1219_p2;
  reg [63:0] xor_ln7_reg_1795;
  wire [63:0] bitcast_ln7_1_fu_1225_p1;
  wire ap_CS_fsm_state70;
  reg [63:0] temp_reg_1805;
  wire ap_CS_fsm_state87;
  wire [3:0] add_ln70_fu_1245_p2;
  reg [3:0] add_ln70_reg_1813;
  wire ap_CS_fsm_state116;
  wire [8:0] add_ln73_1_fu_1295_p2;
  reg [8:0] add_ln73_1_reg_1818;
  wire [0:0] icmp_ln70_fu_1239_p2;
  reg [4:0] deltas_addr_2_reg_1823;
  reg [4:0] activations_addr_6_reg_1828;
  wire [3:0] add_ln72_fu_1307_p2;
  reg [3:0] add_ln72_reg_1836;
  wire ap_CS_fsm_state117;
  wire [0:0] icmp_ln72_fu_1301_p2;
  wire ap_CS_fsm_state128;
  wire [63:0] xor_ln7_2_fu_1346_p2;
  reg [63:0] xor_ln7_2_reg_1856;
  wire ap_CS_fsm_state129;
  wire [63:0] bitcast_ln7_5_fu_1352_p1;
  wire ap_CS_fsm_state130;
  wire [1:0] j_2_fu_1362_p2;
  reg [1:0] j_2_reg_1869;
  wire ap_CS_fsm_state176;
  wire [0:0] icmp_ln123_fu_1356_p2;
  wire [5:0] add_ln90_fu_1392_p2;
  reg [5:0] add_ln90_reg_1874;
  wire [5:0] add_ln90_1_fu_1422_p2;
  reg [5:0] add_ln90_1_reg_1880;
  wire [3:0] select_ln87_fu_1434_p3;
  reg [3:0] select_ln87_reg_1885;
  wire [3:0] ii_1_fu_1447_p2;
  reg [3:0] ii_1_reg_1893;
  wire ap_CS_fsm_state177;
  wire [5:0] add_ln90_2_fu_1457_p2;
  reg [5:0] add_ln90_2_reg_1898;
  wire [0:0] icmp_ln87_fu_1442_p2;
  wire [5:0] add_ln90_4_fu_1467_p2;
  reg [5:0] add_ln90_4_reg_1904;
  wire [8:0] add_ln90_3_fu_1490_p2;
  reg [8:0] add_ln90_3_reg_1915;
  wire [9:0] add_ln90_5_fu_1518_p2;
  reg [9:0] add_ln90_5_reg_1920;
  wire [3:0] jj_2_fu_1530_p2;
  reg [3:0] jj_2_reg_1928;
  wire ap_CS_fsm_state179;
  reg [7:0] weights_addr_2_reg_1933;
  wire [0:0] icmp_ln88_fu_1524_p2;
  reg [8:0] changeMat_addr_1_reg_1943;
  wire [63:0] changeMat_q0;
  reg [63:0] changeMat_load_reg_1948;
  wire ap_CS_fsm_state187;
  reg [4:0] deltas_address0;
  reg deltas_ce0;
  reg deltas_we0;
  reg [63:0] deltas_d0;
  reg [8:0] changeMat_address0;
  reg changeMat_ce0;
  reg changeMat_we0;
  reg [63:0] changeMat_d0;
  reg [4:0] activations_address0;
  reg activations_ce0;
  reg activations_we0;
  reg [63:0] activations_d0;
  reg [1:0] ee_0_reg_324;
  reg [3:0] rows_0_reg_335;
  wire [0:0] icmp_ln159_fu_726_p2;
  reg [3:0] cols_0_reg_346;
  reg [6:0] ee_1_reg_357;
  wire [0:0] icmp_ln167_fu_764_p2;
  reg [6:0] jj_0_reg_368;
  wire [0:0] icmp_ln165_fu_752_p2;
  reg [1:0] cols_1_reg_380;
  wire [0:0] icmp_ln169_fu_860_p2;
  reg [3:0] rows_1_reg_391;
  reg [2:0] i_0_i_reg_402;
  wire ap_CS_fsm_state10;
  reg [1:0] i_1_i_reg_414;
  reg [3:0] ii_0_i_i_reg_425;
  wire ap_CS_fsm_state65;
  reg [3:0] jj_0_i_i_reg_436;
  reg [63:0] x_assign_1_reg_447;
  reg [1:0] i_0_i13_reg_459;
  wire [0:0] icmp_ln111_fu_1148_p2;
  reg [3:0] j_0_i_reg_470;
  reg [3:0] i_0_i_i_reg_481;
  wire ap_CS_fsm_state115;
  reg [3:0] jj_0_i_i21_0_reg_492;
  wire ap_CS_fsm_state175;
  reg [3:0] kk_0_i_i_0_reg_503;
  reg [63:0] error_0_i_i_0_reg_514;
  reg [1:0] level_assign_reg_526;
  reg [3:0] ii_0_i_i25_reg_537;
  reg [3:0] jj_0_i10_i_reg_548;
  wire ap_CS_fsm_state201;
  wire [63:0] zext_ln160_3_fu_691_p1;
  wire [63:0] zext_ln160_7_fu_747_p1;
  wire [63:0] zext_ln170_3_fu_881_p1;
  wire [63:0] zext_ln35_2_fu_907_p1;
  wire [63:0] zext_ln35_fu_912_p1;
  wire [63:0] zext_ln23_4_fu_1026_p1;
  wire [63:0] zext_ln21_5_fu_1087_p1;
  wire [63:0] zext_ln21_3_fu_1051_p1;
  wire [63:0] zext_ln112_3_fu_1169_p1;
  wire [63:0] zext_ln52_5_fu_1199_p1;
  wire [63:0] zext_ln52_6_fu_1210_p1;
  wire [63:0] zext_ln53_fu_1234_p1;
  wire [63:0] zext_ln73_fu_1251_p1;
  wire [63:0] zext_ln73_2_fu_1266_p1;
  wire [63:0] zext_ln73_7_fu_1326_p1;
  wire [63:0] zext_ln73_8_fu_1337_p1;
  wire [63:0] zext_ln90_5_fu_1462_p1;
  wire [63:0] zext_ln90_12_fu_1553_p1;
  wire [63:0] zext_ln89_fu_1563_p1;
  wire [63:0] zext_ln90_13_fu_1573_p1;
  wire ap_CS_fsm_state186;
  wire ap_CS_fsm_state189;
  reg [63:0] grp_fu_559_p0;
  reg [63:0] grp_fu_559_p1;
  wire ap_CS_fsm_state20;
  wire ap_CS_fsm_state38;
  wire ap_CS_fsm_state83;
  wire ap_CS_fsm_state124;
  wire ap_CS_fsm_state143;
  wire ap_CS_fsm_state191;
  wire ap_CS_fsm_state196;
  reg [63:0] grp_fu_566_p0;
  reg [63:0] grp_fu_566_p1;
  wire ap_CS_fsm_state15;
  wire ap_CS_fsm_state110;
  wire ap_CS_fsm_state119;
  wire ap_CS_fsm_state170;
  wire ap_CS_fsm_state181;
  reg [63:0] grp_fu_573_p1;
  wire ap_CS_fsm_state43;
  wire ap_CS_fsm_state88;
  wire ap_CS_fsm_state148;
  reg [63:0] grp_fu_578_p1;
  wire [4:0] tmp_fu_640_p3;
  wire [2:0] tmp_19_fu_652_p3;
  wire [5:0] zext_ln160_1_fu_660_p1;
  wire [5:0] zext_ln160_fu_648_p1;
  wire [5:0] zext_ln160_2_fu_682_p1;
  wire [5:0] add_ln160_1_fu_686_p2;
  wire [8:0] tmp_20_fu_696_p3;
  wire [6:0] tmp_21_fu_708_p3;
  wire [9:0] zext_ln160_4_fu_704_p1;
  wire [9:0] zext_ln160_5_fu_716_p1;
  wire [9:0] zext_ln160_6_fu_738_p1;
  wire [9:0] add_ln160_3_fu_742_p2;
  wire [4:0] tmp_25_fu_788_p3;
  wire [2:0] tmp_26_fu_800_p3;
  wire [5:0] zext_ln170_1_fu_808_p1;
  wire [5:0] zext_ln170_fu_796_p1;
  wire [8:0] tmp_22_fu_818_p3;
  wire [9:0] tmp_23_fu_830_p3;
  wire [7:0] tmp_24_fu_842_p3;
  wire [10:0] zext_ln52_2_fu_850_p1;
  wire [10:0] zext_ln52_1_fu_838_p1;
  wire [5:0] zext_ln170_2_fu_872_p1;
  wire [5:0] add_ln170_1_fu_876_p2;
  wire [9:0] zext_ln35_1_fu_898_p1;
  wire [9:0] add_ln35_fu_902_p2;
  wire [4:0] tmp_27_fu_929_p3;
  wire [2:0] tmp_28_fu_941_p3;
  wire [5:0] zext_ln21_fu_937_p1;
  wire [5:0] zext_ln21_1_fu_949_p1;
  wire [0:0] trunc_ln40_fu_959_p1;
  wire [4:0] tmp_29_fu_971_p3;
  wire [2:0] tmp_30_fu_983_p3;
  wire [5:0] zext_ln23_fu_979_p1;
  wire [5:0] zext_ln23_1_fu_991_p1;
  wire [5:0] zext_ln23_3_fu_1017_p1;
  wire [5:0] add_ln23_1_fu_1021_p2;
  wire [5:0] zext_ln21_2_fu_1042_p1;
  wire [5:0] add_ln21_1_fu_1046_p2;
  wire [6:0] tmp_33_fu_1064_p3;
  wire [8:0] p_shl_cast_fu_1056_p3;
  wire [8:0] zext_ln21_4_fu_1072_p1;
  wire [8:0] add_ln21_2_fu_1076_p2;
  wire [8:0] add_ln21_3_fu_1082_p2;
  wire [63:0] bitcast_ln7_2_fu_1092_p1;
  wire [4:0] tmp_31_fu_1118_p3;
  wire [2:0] tmp_32_fu_1130_p3;
  wire [5:0] zext_ln112_1_fu_1138_p1;
  wire [5:0] zext_ln112_fu_1126_p1;
  wire [5:0] zext_ln112_2_fu_1160_p1;
  wire [5:0] add_ln112_1_fu_1164_p2;
  wire [10:0] zext_ln52_4_fu_1190_p1;
  wire [10:0] add_ln52_1_fu_1194_p2;
  wire [4:0] add_ln52_2_fu_1204_p2;
  wire [63:0] bitcast_ln7_fu_1215_p1;
  wire [4:0] add_ln53_fu_1229_p2;
  wire [4:0] zext_ln73_1_fu_1256_p1;
  wire [4:0] add_ln73_fu_1260_p2;
  wire [7:0] tmp_34_fu_1271_p3;
  wire [5:0] tmp_35_fu_1283_p3;
  wire [8:0] zext_ln73_3_fu_1279_p1;
  wire [8:0] zext_ln73_4_fu_1291_p1;
  wire [8:0] zext_ln73_6_fu_1317_p1;
  wire [8:0] add_ln73_2_fu_1321_p2;
  wire [4:0] zext_ln73_5_fu_1313_p1;
  wire [4:0] add_ln73_3_fu_1331_p2;
  wire [63:0] bitcast_ln7_4_fu_1342_p1;
  wire [4:0] tmp_36_fu_1368_p3;
  wire [2:0] tmp_37_fu_1380_p3;
  wire [5:0] zext_ln90_1_fu_1388_p1;
  wire [5:0] zext_ln90_fu_1376_p1;
  wire [4:0] tmp_38_fu_1398_p3;
  wire [2:0] tmp_39_fu_1410_p3;
  wire [5:0] zext_ln90_3_fu_1418_p1;
  wire [5:0] zext_ln90_2_fu_1406_p1;
  wire [0:0] icmp_ln87_1_fu_1428_p2;
  wire [5:0] zext_ln90_4_fu_1453_p1;
  wire [6:0] tmp_40_fu_1479_p3;
  wire [8:0] p_shl6_cast_fu_1472_p3;
  wire [8:0] zext_ln90_6_fu_1486_p1;
  wire [8:0] tmp_41_fu_1496_p3;
  wire [6:0] tmp_42_fu_1507_p3;
  wire [9:0] zext_ln90_7_fu_1503_p1;
  wire [9:0] zext_ln90_8_fu_1514_p1;
  wire [8:0] zext_ln90_11_fu_1544_p1;
  wire [8:0] add_ln90_6_fu_1548_p2;
  wire [5:0] zext_ln90_10_fu_1540_p1;
  wire [5:0] add_ln89_fu_1558_p2;
  wire [9:0] zext_ln90_9_fu_1536_p1;
  wire [9:0] add_ln90_7_fu_1568_p2;
  reg [1:0] grp_fu_559_opcode;
  reg [200:0] ap_NS_fsm;
  wire Const_0;
  wire Const_1;
  wire [63:0] Const_2;
  wire Const_3;
  wire [63:0] Const_4;
  wire Const_5;
  wire Const_6;
  wire Const_7;
  wire Const_8;
  wire Const_9;
  wire [3:0] Const_10;
  wire Const_11;
  wire Const_12;
  wire Const_13;
  wire Const_14;
  wire [1:0] Const_15;
  wire Const_16;
  wire Const_17;
  wire Const_18;
  wire Const_19;
  wire [1:0] Const_20;
  wire Const_21;
  wire Const_22;
  wire [6:0] Const_23;
  wire Const_24;
  wire Const_25;
  wire Const_26;
  wire Const_27;
  wire Const_28;
  wire [63:0] Const_29;
  wire Const_30;
  wire Const_31;
  wire [1:0] Const_32;
  wire Const_33;
  wire Const_34;
  wire Const_35;
  wire Const_36;
  wire [3:0] Const_37;
  wire Const_38;
  wire Const_39;
  wire Const_40;
  wire Const_41;
  wire [2:0] Const_42;
  wire Const_43;
  wire Const_44;
  wire [1:0] Const_45;
  wire Const_46;
  wire Const_47;
  wire Const_48;
  wire Const_49;
  wire Const_50;
  wire Const_51;
  wire [3:0] Const_52;
  wire Const_53;
  wire Const_54;
  wire Const_55;
  wire [3:0] Const_56;
  wire Const_57;
  wire Const_58;
  wire Const_59;
  wire Const_60;
  wire [3:0] Const_61;
  wire Const_62;
  wire Const_63;
  wire [3:0] Const_64;
  wire Const_65;
  wire Const_66;
  wire Const_67;
  wire [3:0] Const_68;
  wire Const_69;
  wire Const_70;
  wire Const_71;
  wire [3:0] Const_72;
  wire Const_73;
  wire Const_74;
  wire Const_75;
  wire Const_76;
  wire [6:0] Const_77;
  wire Const_78;
  wire Const_79;
  wire Const_80;
  wire [3:0] Const_81;
  wire Const_82;
  wire Const_83;
  wire [1:0] Const_84;
  wire Const_85;
  wire Const_86;
  wire Const_87;
  wire Const_88;
  wire Const_89;
  wire Const_90;
  wire [3:0] Const_91;
  wire Const_92;
  wire Const_93;
  wire Const_94;
  wire Const_95;
  wire [3:0] Const_96;
  wire Const_97;
  wire Const_98;
  wire Const_99;
  wire [63:0] Const_100;
  wire Const_101;
  wire Const_102;
  wire Const_103;
  wire Const_104;
  wire Const_105;
  wire Const_106;
  wire Const_107;
  wire Const_108;
  wire Const_109;
  wire Const_110;
  wire Const_111;
  wire Const_112;
  wire Const_113;
  wire Const_114;
  wire Const_115;
  wire Const_116;
  wire Const_117;
  wire Const_118;
  wire Const_119;
  wire Const_120;
  wire Const_121;
  wire Const_122;
  wire Const_123;
  wire Const_124;
  wire Const_125;
  wire Const_126;
  wire Const_127;
  wire Const_128;
  wire Const_129;
  wire Const_130;
  wire Const_131;
  wire Const_132;
  wire Const_133;
  wire Const_134;
  wire Const_135;
  wire Const_136;
  wire Const_137;
  wire Const_138;
  wire Const_139;
  wire Const_140;
  wire Const_141;
  wire Const_142;
  wire Const_143;
  wire Const_144;
  wire Const_145;
  wire Const_146;
  wire Const_147;
  wire Const_148;
  wire Const_149;
  wire Const_150;
  wire Const_151;
  wire Const_152;
  wire Const_153;
  wire Const_154;
  wire Const_155;
  wire Const_156;
  wire Const_157;
  wire Const_158;
  wire Const_159;
  wire Const_160;
  wire Const_161;
  wire Const_162;
  wire Const_163;
  wire Const_164;
  wire Const_165;
  wire Const_166;
  wire Const_167;
  wire Const_168;
  wire Const_169;
  wire Const_170;
  wire Const_171;
  wire Const_172;
  wire Const_173;
  wire Const_174;
  wire Const_175;
  wire Const_176;
  wire Const_177;
  wire Const_178;
  wire Const_179;
  wire Const_180;
  wire Const_181;
  wire Const_182;
  wire Const_183;
  wire Const_184;
  wire Const_185;
  wire Const_186;
  wire Const_187;
  wire Const_188;
  wire Const_189;
  wire Const_190;
  wire Const_191;
  wire Const_192;
  wire Const_193;
  wire Const_194;
  wire [63:0] Const_195;
  wire Const_196;
  wire Const_197;
  wire Const_198;
  wire Const_199;
  wire Const_200;
  wire Const_201;
  wire Const_202;
  wire Const_203;
  wire Const_204;
  wire Const_205;
  wire Const_206;
  wire Const_207;
  wire Const_208;
  wire Const_209;
  wire Const_210;
  wire Const_211;
  wire Const_212;
  wire Const_213;
  wire Const_214;
  wire Const_215;
  wire Const_216;
  wire Const_217;
  wire Const_218;
  wire Const_219;
  wire Const_220;
  wire Const_221;
  wire Const_222;
  wire Const_223;
  wire [63:0] Const_224;
  wire Const_225;
  wire Const_226;
  wire Const_227;
  wire Const_228;
  wire Const_229;
  wire Const_230;
  wire Const_231;
  wire Const_232;
  wire Const_233;
  wire Const_234;
  wire Const_235;
  wire Const_236;
  wire Const_237;
  wire Const_238;
  wire Const_239;
  wire Const_240;
  wire Const_241;
  wire Const_242;
  wire Const_243;
  wire Const_244;
  wire [63:0] Const_245;
  wire Const_246;
  wire Const_247;
  wire Const_248;
  wire Const_249;
  wire Const_250;
  wire Const_251;
  wire Const_252;
  wire [1:0] Const_253;
  wire Const_254;
  wire Const_255;
  wire Const_256;
  wire Const_257;
  wire Const_258;
  wire Const_259;
  wire Const_260;
  wire [1:0] Const_261;
  wire Const_262;
  wire Const_263;
  wire Const_264;
  wire Const_265;
  wire Const_266;
  wire Const_267;
  wire Const_268;
  wire Const_269;
  wire Const_270;
  wire Const_271;
  wire Const_272;
  wire Const_273;
  wire [63:0] Const_274;
  wire Const_275;
  wire Const_276;
  wire Const_277;
  wire Const_278;
  wire Const_279;
  wire Const_280;
  wire Const_281;
  wire Const_282;
  wire Const_283;
  wire Const_284;
  wire Const_285;
  wire Const_286;
  wire [63:0] Const_287;
  wire Const_288;
  wire [63:0] Const_289;
  wire Const_290;
  wire Const_291;
  wire Const_292;
  wire Const_293;
  wire Const_294;
  wire Const_295;
  wire Const_296;
  wire Const_297;
  wire Const_298;
  wire Const_299;
  wire Const_300;
  wire Const_301;
  wire Const_302;
  wire Const_303;
  wire Const_304;
  wire Const_305;
  wire Const_306;
  wire Const_307;
  wire Const_308;
  wire Const_309;
  wire Const_310;
  wire Const_311;
  wire Const_312;
  wire Const_313;
  wire Const_314;
  wire Const_315;
  wire Const_316;
  wire Const_317;
  wire Const_318;
  wire Const_319;
  wire Const_320;
  wire Const_321;
  wire Const_322;
  wire Const_323;
  wire Const_324;
  wire Const_325;
  wire Const_326;
  wire Const_327;
  wire Const_328;
  wire Const_329;
  wire Const_330;
  wire Const_331;
  wire Const_332;
  wire Const_333;
  wire Const_334;
  wire Const_335;
  wire Const_336;
  wire Const_337;
  wire Const_338;
  wire Const_339;
  wire Const_340;
  wire Const_341;
  wire Const_342;
  wire Const_343;
  wire Const_344;
  wire Const_345;
  wire Const_346;
  wire Const_347;
  wire Const_348;
  wire Const_349;
  wire Const_350;
  wire Const_351;
  wire Const_352;
  wire Const_353;
  wire Const_354;
  wire Const_355;
  wire Const_356;
  wire Const_357;
  wire Const_358;
  wire Const_359;
  wire [4:0] Const_360;
  wire [4:0] Const_361;
  wire [3:0] Const_362;
  wire [3:0] Const_363;
  wire [4:0] Const_364;
  wire [4:0] Const_365;
  wire [1:0] Const_366;
  wire [3:0] Const_367;
  wire [6:0] Const_368;
  wire [1:0] Const_369;
  wire [1:0] Const_370;
  wire [3:0] Const_371;
  wire [1:0] Const_372;
  wire [2:0] Const_373;
  wire [1:0] Const_374;
  wire Const_375;
  wire Const_376;
  wire [3:0] Const_377;
  wire Const_378;
  wire Const_379;
  wire [1:0] Const_380;
  wire Const_381;
  wire Const_382;
  wire [1:0] Const_383;
  wire Const_384;
  wire Const_385;
  wire [3:0] Const_386;
  wire Const_387;
  wire Const_388;
  wire [3:0] Const_389;
  wire Const_390;
  wire Const_391;
  wire [6:0] Const_392;
  wire Const_393;
  wire Const_394;
  wire [6:0] Const_395;
  wire Const_396;
  wire Const_397;
  wire [1:0] Const_398;
  wire Const_399;
  wire Const_400;
  wire [3:0] Const_401;
  wire Const_402;
  wire Const_403;
  wire [3:0] Const_404;
  wire Const_405;
  wire Const_406;
  wire Const_407;
  wire Const_408;
  wire [2:0] Const_409;
  wire Const_410;
  wire Const_411;
  wire [1:0] Const_412;
  wire Const_413;
  wire Const_414;
  wire [3:0] Const_415;
  wire Const_416;
  wire Const_417;
  wire [3:0] Const_418;
  wire Const_419;
  wire Const_420;
  wire [3:0] Const_421;
  wire Const_422;
  wire Const_423;
  wire [1:0] Const_424;
  wire Const_425;
  wire Const_426;
  wire Const_427;
  wire Const_428;
  wire [3:0] Const_429;
  wire Const_430;
  wire Const_431;
  wire [3:0] Const_432;
  wire [3:0] Const_433;
  wire [1:0] Const_434;
  wire [3:0] Const_435;
  wire [6:0] Const_436;
  wire [3:0] Const_437;
  wire [3:0] Const_438;
  wire [3:0] Const_439;
  wire [3:0] Const_440;
  wire Const_441;
  wire [3:0] Const_442;
  wire [3:0] Const_443;
  wire Const_444;
  wire [3:0] Const_445;
  wire [3:0] Const_446;
  wire [63:0] Const_447;
  wire [63:0] Const_448;
  wire [63:0] Const_449;
  input [3070:0] locking_key;
  wire [1653:0] working_key;

  initial begin
    #0 ap_CS_fsm = 201'd1;
  end


  backprop_deltas
  #(
    .DataWidth(64),
    .AddressRange(30),
    .AddressWidth(5)
  )
  deltas_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(deltas_address0),
    .ce0(deltas_ce0),
    .we0(deltas_we0),
    .d0(deltas_d0),
    .q0(deltas_q0)
  );


  backprop_changeMat
  #(
    .DataWidth(64),
    .AddressRange(300),
    .AddressWidth(9)
  )
  changeMat_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(changeMat_address0),
    .ce0(changeMat_ce0),
    .we0(changeMat_we0),
    .d0(changeMat_d0),
    .q0(changeMat_q0)
  );


  backprop_deltas
  #(
    .DataWidth(64),
    .AddressRange(30),
    .AddressWidth(5)
  )
  activations_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(activations_address0),
    .ce0(activations_ce0),
    .we0(activations_we0),
    .d0(activations_d0),
    .q0(activations_q0)
  );

  assign Const_0 = (1'd1 ^ working_key[0]);

  backprop_dadddsubcud
  #(
    .ID(1),
    .NUM_STAGE(5),
    .din0_WIDTH(64),
    .din1_WIDTH(64),
    .dout_WIDTH(64)
  )
  backprop_dadddsubcud_U1
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_559_p0),
    .din1(grp_fu_559_p1),
    .opcode(grp_fu_559_opcode),
    .ce(Const_0),
    .dout(grp_fu_559_p2)
  );

  assign Const_1 = (1'd0 ^ working_key[1]);

  backprop_dmul_64ndEe
  #(
    .ID(1),
    .NUM_STAGE(5),
    .din0_WIDTH(64),
    .din1_WIDTH(64),
    .dout_WIDTH(64)
  )
  backprop_dmul_64ndEe_U2
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_566_p0),
    .din1(grp_fu_566_p1),
    .ce(Const_1),
    .dout(grp_fu_566_p2)
  );

  assign Const_2 = (64'd15445740152669152618 ^ working_key[65:2]);
  assign Const_3 = (1'd0 ^ working_key[66]);

  backprop_ddiv_64neOg
  #(
    .ID(1),
    .NUM_STAGE(22),
    .din0_WIDTH(64),
    .din1_WIDTH(64),
    .dout_WIDTH(64)
  )
  backprop_ddiv_64neOg_U3
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(Const_2),
    .din1(grp_fu_573_p1),
    .ce(Const_3),
    .dout(grp_fu_573_p2)
  );

  assign Const_4 = (64'd5524415532170389847 ^ working_key[130:67]);
  assign Const_5 = (1'd0 ^ working_key[131]);

  backprop_dexp_64nfYi
  #(
    .ID(1),
    .NUM_STAGE(13),
    .din0_WIDTH(64),
    .din1_WIDTH(64),
    .dout_WIDTH(64)
  )
  backprop_dexp_64nfYi_U4
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(Const_4),
    .din1(grp_fu_578_p1),
    .ce(Const_5),
    .dout(grp_fu_578_p2)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end

  assign Const_6 = (1'd0 ^ working_key[132]);
  assign Const_7 = (1'd0 ^ working_key[133]);
  assign Const_8 = (1'd0 ^ working_key[134]);
  assign Const_9 = (1'd0 ^ working_key[135]);
  assign Const_10 = (4'd5 ^ working_key[139:136]);

  always @(posedge ap_clk) begin
    if(((icmp_ln159_fu_726_p2 == Const_6) & (Const_7 == ap_CS_fsm_state4) ^ working_key[140]) == 1'b0) begin
      cols_0_reg_346 <= cols_fu_732_p2;
    end else if((icmp_ln157_fu_670_p2 == Const_8) & (Const_9 == ap_CS_fsm_state3)) begin
      cols_0_reg_346 <= Const_10;
    end 
  end

  assign Const_11 = (1'd1 ^ working_key[141]);
  assign Const_12 = (1'd1 ^ working_key[142]);
  assign Const_13 = (1'd1 ^ working_key[143]);
  assign Const_14 = (1'd1 ^ working_key[144]);
  assign Const_15 = (2'd2 ^ working_key[146:145]);

  always @(posedge ap_clk) begin
    if(((icmp_ln169_fu_860_p2 == Const_11) & (Const_12 == ap_CS_fsm_state8) ^ working_key[147]) == 1'b1) begin
      cols_1_reg_380 <= cols_2_reg_1631;
    end else if((icmp_ln167_fu_764_p2 == Const_13) & (Const_14 == ap_CS_fsm_state6)) begin
      cols_1_reg_380 <= Const_15;
    end 
  end

  assign Const_16 = (1'd0 ^ working_key[148]);
  assign Const_17 = (1'd1 ^ working_key[149]);
  assign Const_18 = (1'd0 ^ working_key[150]);
  assign Const_19 = (1'd1 ^ working_key[151]);
  assign Const_20 = (2'd3 ^ working_key[153:152]);

  always @(posedge ap_clk) begin
    if(((icmp_ln157_fu_670_p2 == Const_16) & (Const_17 == ap_CS_fsm_state3) ^ working_key[154]) == 1'b1) begin
      ee_0_reg_324 <= ee_reg_1581;
    end else if((ap_start == Const_18) & (Const_19 == ap_CS_fsm_state1)) begin
      ee_0_reg_324 <= Const_20;
    end 
  end

  assign Const_21 = (1'd1 ^ working_key[155]);
  assign Const_22 = (1'd0 ^ working_key[156]);
  assign Const_23 = (7'd46 ^ working_key[163:157]);
  assign Const_24 = (1'd0 ^ working_key[164]);
  assign Const_25 = (1'd1 ^ working_key[165]);

  always @(posedge ap_clk) begin
    if(((icmp_ln156_fu_628_p2 == Const_21) & (Const_22 == ap_CS_fsm_state2) ^ working_key[166]) == 1'b0) begin
      ee_1_reg_357 <= Const_23;
    end else if((icmp_ln167_fu_764_p2 == Const_24) & (Const_25 == ap_CS_fsm_state6)) begin
      ee_1_reg_357 <= ee_2_reg_1615;
    end 
  end

  assign Const_26 = (1'd1 ^ working_key[167]);
  assign Const_27 = (1'd1 ^ working_key[168]);
  assign Const_28 = (1'd0 ^ working_key[169]);
  assign Const_29 = (64'd5788626709681646154 ^ working_key[233:170]);

  always @(posedge ap_clk) begin
    if(((Const_26 == ap_CS_fsm_state128) ^ working_key[234]) == 1'b0) begin
      error_0_i_i_0_reg_514 <= grp_fu_559_p2;
    end else if((icmp_ln70_fu_1239_p2 == Const_27) & (Const_28 == ap_CS_fsm_state116)) begin
      error_0_i_i_0_reg_514 <= Const_29;
    end 
  end

  assign Const_30 = (1'd1 ^ working_key[235]);
  assign Const_31 = (1'd0 ^ working_key[236]);
  assign Const_32 = (2'd2 ^ working_key[238:237]);
  assign Const_33 = (1'd1 ^ working_key[239]);
  assign Const_34 = (1'd0 ^ working_key[240]);

  always @(posedge ap_clk) begin
    if(((icmp_ln39_fu_917_p2 == Const_30) & (Const_31 == ap_CS_fsm_state11) ^ working_key[241]) == 1'b1) begin
      i_0_i13_reg_459 <= Const_32;
    end else if((icmp_ln111_fu_1148_p2 == Const_33) & (Const_34 == ap_CS_fsm_state67)) begin
      i_0_i13_reg_459 <= i_3_reg_1749;
    end 
  end

  assign Const_35 = (1'd0 ^ working_key[242]);
  assign Const_36 = (1'd1 ^ working_key[243]);
  assign Const_37 = (4'd5 ^ working_key[247:244]);
  assign Const_38 = (1'd0 ^ working_key[248]);

  always @(posedge ap_clk) begin
    if(((icmp_ln110_fu_1106_p2 == Const_35) & (Const_36 == ap_CS_fsm_state66) ^ working_key[249]) == 1'b1) begin
      i_0_i_i_reg_481 <= Const_37;
    end else if(Const_38 == ap_CS_fsm_state115) begin
      i_0_i_i_reg_481 <= i_2_reg_1770;
    end 
  end

  assign Const_39 = (1'd0 ^ working_key[250]);
  assign Const_40 = (1'd1 ^ working_key[251]);
  assign Const_41 = (1'd1 ^ working_key[252]);
  assign Const_42 = (3'd3 ^ working_key[255:253]);

  always @(posedge ap_clk) begin
    if(((Const_39 == ap_CS_fsm_state10) ^ working_key[256]) == 1'b0) begin
      i_0_i_reg_402 <= i_reg_1662;
    end else if((icmp_ln168_fu_776_p2 == Const_40) & (Const_41 == ap_CS_fsm_state7)) begin
      i_0_i_reg_402 <= Const_42;
    end 
  end

  assign Const_43 = (1'd0 ^ working_key[257]);
  assign Const_44 = (1'd0 ^ working_key[258]);
  assign Const_45 = (2'd1 ^ working_key[260:259]);
  assign Const_46 = (1'd0 ^ working_key[261]);
  assign Const_47 = (1'd1 ^ working_key[262]);

  always @(posedge ap_clk) begin
    if(((icmp_ln34_fu_886_p2 == Const_43) & (Const_44 == ap_CS_fsm_state9) ^ working_key[263]) == 1'b0) begin
      i_1_i_reg_414 <= Const_45;
    end else if((icmp_ln18_fu_1001_p2 == Const_46) & (Const_47 == ap_CS_fsm_state12)) begin
      i_1_i_reg_414 <= i_1_reg_1675;
    end 
  end

  assign Const_48 = (1'd0 ^ working_key[264]);
  assign Const_49 = (1'd1 ^ working_key[265]);
  assign Const_50 = (1'd1 ^ working_key[266]);
  assign Const_51 = (1'd1 ^ working_key[267]);
  assign Const_52 = (4'd9 ^ working_key[271:268]);

  always @(posedge ap_clk) begin
    if(((icmp_ln88_fu_1524_p2 == Const_48) & (Const_49 == ap_CS_fsm_state179) ^ working_key[272]) == 1'b1) begin
      ii_0_i_i25_reg_537 <= ii_1_reg_1893;
    end else if((icmp_ln123_fu_1356_p2 == Const_50) & (Const_51 == ap_CS_fsm_state176)) begin
      ii_0_i_i25_reg_537 <= Const_52;
    end 
  end

  assign Const_53 = (1'd1 ^ working_key[273]);
  assign Const_54 = (1'd1 ^ working_key[274]);
  assign Const_55 = (1'd1 ^ working_key[275]);
  assign Const_56 = (4'd5 ^ working_key[279:276]);

  always @(posedge ap_clk) begin
    if(((Const_53 == ap_CS_fsm_state65) ^ working_key[280]) == 1'b0) begin
      ii_0_i_i_reg_425 <= ii_reg_1698;
    end else if((icmp_ln39_fu_917_p2 == Const_54) & (Const_55 == ap_CS_fsm_state11)) begin
      ii_0_i_i_reg_425 <= Const_56;
    end 
  end

  assign Const_57 = (1'd1 ^ working_key[281]);
  assign Const_58 = (1'd1 ^ working_key[282]);
  assign Const_59 = (1'd0 ^ working_key[283]);
  assign Const_60 = (1'd0 ^ working_key[284]);
  assign Const_61 = (4'd14 ^ working_key[288:285]);

  always @(posedge ap_clk) begin
    if(((icmp_ln111_fu_1148_p2 == Const_57) & (Const_58 == ap_CS_fsm_state67) ^ working_key[289]) == 1'b1) begin
      j_0_i_reg_470 <= j_fu_1154_p2;
    end else if((icmp_ln110_fu_1106_p2 == Const_59) & (Const_60 == ap_CS_fsm_state66)) begin
      j_0_i_reg_470 <= Const_61;
    end 
  end

  assign Const_62 = (1'd0 ^ working_key[290]);
  assign Const_63 = (1'd1 ^ working_key[291]);
  assign Const_64 = (4'd5 ^ working_key[295:292]);

  always @(posedge ap_clk) begin
    if(((Const_62 == ap_CS_fsm_state201) ^ working_key[296]) == 1'b0) begin
      jj_0_i10_i_reg_548 <= jj_2_reg_1928;
    end else if(Const_63 == ap_CS_fsm_state178) begin
      jj_0_i10_i_reg_548 <= Const_64;
    end 
  end

  assign Const_65 = (1'd0 ^ working_key[297]);
  assign Const_66 = (1'd1 ^ working_key[298]);
  assign Const_67 = (1'd0 ^ working_key[299]);
  assign Const_68 = (4'd2 ^ working_key[303:300]);

  always @(posedge ap_clk) begin
    if(((Const_65 == ap_CS_fsm_state175) ^ working_key[304]) == 1'b0) begin
      jj_0_i_i21_0_reg_492 <= add_ln70_reg_1813;
    end else if((icmp_ln51_fu_1174_p2 == Const_66) & (Const_67 == ap_CS_fsm_state68)) begin
      jj_0_i_i21_0_reg_492 <= Const_68;
    end 
  end

  assign Const_69 = (1'd1 ^ working_key[305]);
  assign Const_70 = (1'd0 ^ working_key[306]);
  assign Const_71 = (1'd0 ^ working_key[307]);
  assign Const_72 = (4'd10 ^ working_key[311:308]);

  always @(posedge ap_clk) begin
    if(((Const_69 == ap_CS_fsm_state24) ^ working_key[312]) == 1'b1) begin
      jj_0_i_i_reg_436 <= jj_reg_1716;
    end else if((icmp_ln18_fu_1001_p2 == Const_70) & (Const_71 == ap_CS_fsm_state12)) begin
      jj_0_i_i_reg_436 <= Const_72;
    end 
  end

  assign Const_73 = (1'd0 ^ working_key[313]);
  assign Const_74 = (1'd0 ^ working_key[314]);
  assign Const_75 = (1'd0 ^ working_key[315]);
  assign Const_76 = (1'd1 ^ working_key[316]);
  assign Const_77 = (7'd125 ^ working_key[323:317]);

  always @(posedge ap_clk) begin
    if(((icmp_ln123_fu_1356_p2 == Const_73) & (Const_74 == ap_CS_fsm_state176) ^ working_key[324]) == 1'b0) begin
      jj_0_reg_368 <= jj_1_reg_1623;
    end else if((icmp_ln165_fu_752_p2 == Const_75) & (Const_76 == ap_CS_fsm_state5)) begin
      jj_0_reg_368 <= Const_77;
    end 
  end

  assign Const_78 = (1'd0 ^ working_key[325]);
  assign Const_79 = (1'd0 ^ working_key[326]);
  assign Const_80 = (1'd0 ^ working_key[327]);
  assign Const_81 = (4'd10 ^ working_key[331:328]);

  always @(posedge ap_clk) begin
    if(((Const_78 == ap_CS_fsm_state128) ^ working_key[332]) == 1'b1) begin
      kk_0_i_i_0_reg_503 <= add_ln72_reg_1836;
    end else if((icmp_ln70_fu_1239_p2 == Const_79) & (Const_80 == ap_CS_fsm_state116)) begin
      kk_0_i_i_0_reg_503 <= Const_81;
    end 
  end

  assign Const_82 = (1'd1 ^ working_key[333]);
  assign Const_83 = (1'd0 ^ working_key[334]);
  assign Const_84 = (2'd0 ^ working_key[336:335]);
  assign Const_85 = (1'd0 ^ working_key[337]);
  assign Const_86 = (1'd0 ^ working_key[338]);

  always @(posedge ap_clk) begin
    if(((icmp_ln70_fu_1239_p2 == Const_82) & (Const_83 == ap_CS_fsm_state116) ^ working_key[339]) == 1'b1) begin
      level_assign_reg_526 <= Const_84;
    end else if((icmp_ln87_fu_1442_p2 == Const_85) & (Const_86 == ap_CS_fsm_state177)) begin
      level_assign_reg_526 <= j_2_reg_1869;
    end 
  end

  assign Const_87 = (1'd0 ^ working_key[340]);
  assign Const_88 = (1'd1 ^ working_key[341]);
  assign Const_89 = (1'd1 ^ working_key[342]);
  assign Const_90 = (1'd1 ^ working_key[343]);
  assign Const_91 = (4'd5 ^ working_key[347:344]);

  always @(posedge ap_clk) begin
    if(((icmp_ln159_fu_726_p2 == Const_87) & (Const_88 == ap_CS_fsm_state4) ^ working_key[348]) == 1'b0) begin
      rows_0_reg_335 <= rows_reg_1594;
    end else if((icmp_ln156_fu_628_p2 == Const_89) & (Const_90 == ap_CS_fsm_state2)) begin
      rows_0_reg_335 <= Const_91;
    end 
  end

  assign Const_92 = (1'd0 ^ working_key[349]);
  assign Const_93 = (1'd0 ^ working_key[350]);
  assign Const_94 = (1'd0 ^ working_key[351]);
  assign Const_95 = (1'd0 ^ working_key[352]);
  assign Const_96 = (4'd0 ^ working_key[356:353]);

  always @(posedge ap_clk) begin
    if(((icmp_ln169_fu_860_p2 == Const_92) & (Const_93 == ap_CS_fsm_state8) ^ working_key[357]) == 1'b1) begin
      rows_1_reg_391 <= rows_2_fu_866_p2;
    end else if((icmp_ln168_fu_776_p2 == Const_94) & (Const_95 == ap_CS_fsm_state7)) begin
      rows_1_reg_391 <= Const_96;
    end 
  end

  assign Const_97 = (1'd0 ^ working_key[358]);
  assign Const_98 = (1'd0 ^ working_key[359]);
  assign Const_99 = (1'd0 ^ working_key[360]);
  assign Const_100 = (64'd12315561894402501290 ^ working_key[424:361]);

  always @(posedge ap_clk) begin
    if(((Const_97 == ap_CS_fsm_state24) ^ working_key[425]) == 1'b0) begin
      x_assign_1_reg_447 <= grp_fu_559_p2;
    end else if((icmp_ln18_fu_1001_p2 == Const_98) & (Const_99 == ap_CS_fsm_state12)) begin
      x_assign_1_reg_447 <= Const_100;
    end 
  end

  assign Const_101 = (1'd0 ^ working_key[426]);
  assign Const_102 = (1'd0 ^ working_key[427]);

  always @(posedge ap_clk) begin
    if((icmp_ln18_fu_1001_p2 == Const_101) & (Const_102 == ap_CS_fsm_state12)) begin
      activations_addr_5_reg_1708 <= zext_ln23_4_fu_1026_p1;
      zext_ln23_2_reg_1703[3:0] <= zext_ln23_2_fu_1013_p1[3:0];
    end 
  end

  assign Const_103 = (1'd0 ^ working_key[428]);
  assign Const_104 = (1'd0 ^ working_key[429]);

  always @(posedge ap_clk) begin
    if((icmp_ln70_fu_1239_p2 == Const_103) & (Const_104 == ap_CS_fsm_state116)) begin
      activations_addr_6_reg_1828 <= zext_ln73_2_fu_1266_p1;
      add_ln73_1_reg_1818[8:1] <= add_ln73_1_fu_1295_p2[8:1];
      deltas_addr_2_reg_1823[3:0] <= zext_ln73_fu_1251_p1[3:0];
    end 
  end

  assign Const_105 = (1'd0 ^ working_key[430]);
  assign Const_106 = (1'd1 ^ working_key[431]);

  always @(posedge ap_clk) begin
    if((icmp_ln110_fu_1106_p2 == Const_105) & (Const_106 == ap_CS_fsm_state66)) begin
      add_ln112_reg_1754[5:1] <= add_ln112_fu_1142_p2[5:1];
    end 
  end

  assign Const_107 = (1'd1 ^ working_key[432]);
  assign Const_108 = (1'd1 ^ working_key[433]);

  always @(posedge ap_clk) begin
    if((icmp_ln157_fu_670_p2 == Const_107) & (Const_108 == ap_CS_fsm_state3)) begin
      add_ln160_2_reg_1599[9:1] <= add_ln160_2_fu_720_p2[9:1];
    end 
  end

  assign Const_109 = (1'd0 ^ working_key[434]);
  assign Const_110 = (1'd0 ^ working_key[435]);

  always @(posedge ap_clk) begin
    if((icmp_ln156_fu_628_p2 == Const_109) & (Const_110 == ap_CS_fsm_state2)) begin
      add_ln160_reg_1586[5:1] <= add_ln160_fu_664_p2[5:1];
    end 
  end

  assign Const_111 = (1'd0 ^ working_key[436]);
  assign Const_112 = (1'd0 ^ working_key[437]);

  always @(posedge ap_clk) begin
    if((icmp_ln168_fu_776_p2 == Const_111) & (Const_112 == ap_CS_fsm_state7)) begin
      add_ln170_reg_1636[5:1] <= add_ln170_fu_812_p2[5:1];
    end 
  end

  assign Const_113 = (1'd0 ^ working_key[438]);
  assign Const_114 = (1'd0 ^ working_key[439]);

  always @(posedge ap_clk) begin
    if((icmp_ln39_fu_917_p2 == Const_113) & (Const_114 == ap_CS_fsm_state11)) begin
      add_ln21_reg_1680[5:1] <= add_ln21_fu_953_p2[5:1];
      add_ln23_reg_1690[5:1] <= add_ln23_fu_995_p2[5:1];
      select_ln40_reg_1685[3:1] <= select_ln40_fu_963_p3[3:1];
    end 
  end

  assign Const_115 = (1'd1 ^ working_key[440]);
  assign Const_116 = (1'd0 ^ working_key[441]);

  always @(posedge ap_clk) begin
    if((icmp_ln168_fu_776_p2 == Const_115) & (Const_116 == ap_CS_fsm_state7)) begin
      add_ln52_reg_1646[10:1] <= add_ln52_fu_854_p2[10:1];
      zext_ln52_reg_1641[8:2] <= zext_ln52_fu_826_p1[8:2];
    end 
  end

  assign Const_117 = (1'd0 ^ working_key[442]);

  always @(posedge ap_clk) begin
    if(Const_117 == ap_CS_fsm_state116) begin
      add_ln70_reg_1813 <= add_ln70_fu_1245_p2;
    end 
  end

  assign Const_118 = (1'd1 ^ working_key[443]);

  always @(posedge ap_clk) begin
    if(Const_118 == ap_CS_fsm_state117) begin
      add_ln72_reg_1836 <= add_ln72_fu_1307_p2;
    end 
  end

  assign Const_119 = (1'd0 ^ working_key[444]);
  assign Const_120 = (1'd0 ^ working_key[445]);

  always @(posedge ap_clk) begin
    if((icmp_ln123_fu_1356_p2 == Const_119) & (Const_120 == ap_CS_fsm_state176)) begin
      add_ln90_1_reg_1880[5:1] <= add_ln90_1_fu_1422_p2[5:1];
      add_ln90_reg_1874[5:1] <= add_ln90_fu_1392_p2[5:1];
      j_2_reg_1869 <= j_2_fu_1362_p2;
      select_ln87_reg_1885[3:1] <= select_ln87_fu_1434_p3[3:1];
    end 
  end

  assign Const_121 = (1'd1 ^ working_key[446]);
  assign Const_122 = (1'd0 ^ working_key[447]);

  always @(posedge ap_clk) begin
    if((icmp_ln87_fu_1442_p2 == Const_121) & (Const_122 == ap_CS_fsm_state177)) begin
      add_ln90_2_reg_1898 <= add_ln90_2_fu_1457_p2;
      add_ln90_4_reg_1904 <= add_ln90_4_fu_1467_p2;
    end 
  end

  assign Const_123 = (1'd0 ^ working_key[448]);

  always @(posedge ap_clk) begin
    if(Const_123 == ap_CS_fsm_state178) begin
      add_ln90_3_reg_1915[8:1] <= add_ln90_3_fu_1490_p2[8:1];
      add_ln90_5_reg_1920[9:1] <= add_ln90_5_fu_1518_p2[9:1];
    end 
  end

  assign Const_124 = (1'd1 ^ working_key[449]);
  assign Const_125 = (1'd0 ^ working_key[450]);

  always @(posedge ap_clk) begin
    if((icmp_ln88_fu_1524_p2 == Const_124) & (Const_125 == ap_CS_fsm_state179)) begin
      changeMat_addr_1_reg_1943 <= zext_ln90_13_fu_1573_p1;
      weights_addr_2_reg_1933 <= zext_ln90_12_fu_1553_p1;
    end 
  end

  assign Const_126 = (1'd0 ^ working_key[451]);

  always @(posedge ap_clk) begin
    if(Const_126 == ap_CS_fsm_state187) begin
      changeMat_load_reg_1948 <= changeMat_q0;
    end 
  end

  assign Const_127 = (1'd0 ^ working_key[452]);

  always @(posedge ap_clk) begin
    if(Const_127 == ap_CS_fsm_state7) begin
      cols_2_reg_1631 <= cols_2_fu_782_p2;
    end 
  end

  assign Const_128 = (1'd0 ^ working_key[453]);

  always @(posedge ap_clk) begin
    if(Const_128 == ap_CS_fsm_state5) begin
      ee_2_reg_1615 <= ee_2_fu_758_p2;
    end 
  end

  assign Const_129 = (1'd1 ^ working_key[454]);

  always @(posedge ap_clk) begin
    if(Const_129 == ap_CS_fsm_state2) begin
      ee_reg_1581 <= ee_fu_634_p2;
    end 
  end

  assign Const_130 = (1'd0 ^ working_key[455]);

  always @(posedge ap_clk) begin
    if(Const_130 == ap_CS_fsm_state11) begin
      i_1_reg_1675 <= i_1_fu_923_p2;
    end 
  end

  assign Const_131 = (1'd1 ^ working_key[456]);

  always @(posedge ap_clk) begin
    if(Const_131 == ap_CS_fsm_state68) begin
      i_2_reg_1770 <= i_2_fu_1180_p2;
    end 
  end

  assign Const_132 = (1'd0 ^ working_key[457]);

  always @(posedge ap_clk) begin
    if(Const_132 == ap_CS_fsm_state66) begin
      i_3_reg_1749 <= i_3_fu_1112_p2;
    end 
  end

  assign Const_133 = (1'd1 ^ working_key[458]);

  always @(posedge ap_clk) begin
    if(Const_133 == ap_CS_fsm_state9) begin
      i_reg_1662 <= i_fu_892_p2;
    end 
  end

  assign Const_134 = (1'd0 ^ working_key[459]);

  always @(posedge ap_clk) begin
    if(Const_134 == ap_CS_fsm_state177) begin
      ii_1_reg_1893 <= ii_1_fu_1447_p2;
    end 
  end

  assign Const_135 = (1'd1 ^ working_key[460]);

  always @(posedge ap_clk) begin
    if(Const_135 == ap_CS_fsm_state12) begin
      ii_reg_1698 <= ii_fu_1007_p2;
    end 
  end

  assign Const_136 = (1'd1 ^ working_key[461]);

  always @(posedge ap_clk) begin
    if(Const_136 == ap_CS_fsm_state6) begin
      jj_1_reg_1623 <= jj_1_fu_770_p2;
    end 
  end

  assign Const_137 = (1'd0 ^ working_key[462]);

  always @(posedge ap_clk) begin
    if(Const_137 == ap_CS_fsm_state179) begin
      jj_2_reg_1928 <= jj_2_fu_1530_p2;
    end 
  end

  assign Const_138 = (1'd1 ^ working_key[463]);

  always @(posedge ap_clk) begin
    if(Const_138 == ap_CS_fsm_state13) begin
      jj_reg_1716 <= jj_fu_1036_p2;
    end 
  end

  assign Const_139 = (1'd0 ^ working_key[464]);
  assign Const_140 = (1'd1 ^ working_key[465]);
  assign Const_141 = (1'd0 ^ working_key[466]);

  always @(posedge ap_clk) begin
    if((Const_139 == ap_CS_fsm_state178) | (Const_140 == ap_CS_fsm_state69) | (Const_141 == ap_CS_fsm_state14)) begin
      reg_583 <= activations_q0;
    end 
  end

  assign Const_142 = (1'd1 ^ working_key[467]);
  assign Const_143 = (1'd0 ^ working_key[468]);
  assign Const_144 = (1'd1 ^ working_key[469]);

  always @(posedge ap_clk) begin
    if((Const_142 == ap_CS_fsm_state190) | (Const_143 == ap_CS_fsm_state118) | (Const_144 == ap_CS_fsm_state14)) begin
      reg_590 <= weights_q0;
    end 
  end

  assign Const_145 = (1'd0 ^ working_key[470]);
  assign Const_146 = (1'd1 ^ working_key[471]);
  assign Const_147 = (1'd0 ^ working_key[472]);
  assign Const_148 = (1'd1 ^ working_key[473]);
  assign Const_149 = (1'd0 ^ working_key[474]);
  assign Const_150 = (1'd1 ^ working_key[475]);
  assign Const_151 = (1'd0 ^ working_key[476]);

  always @(posedge ap_clk) begin
    if((Const_145 == ap_CS_fsm_state195) | (Const_146 == ap_CS_fsm_state185) | (Const_147 == ap_CS_fsm_state174) | (Const_148 == ap_CS_fsm_state123) | (Const_149 == ap_CS_fsm_state114) | (Const_150 == ap_CS_fsm_state19) | (Const_151 == ap_CS_fsm_state190)) begin
      reg_596 <= grp_fu_566_p2;
    end 
  end

  assign Const_152 = (1'd1 ^ working_key[477]);
  assign Const_153 = (1'd0 ^ working_key[478]);
  assign Const_154 = (1'd1 ^ working_key[479]);

  always @(posedge ap_clk) begin
    if((Const_152 == ap_CS_fsm_state142) | (Const_153 == ap_CS_fsm_state82) | (Const_154 == ap_CS_fsm_state37)) begin
      reg_604 <= grp_fu_578_p2;
    end 
  end

  assign Const_155 = (1'd0 ^ working_key[480]);
  assign Const_156 = (1'd1 ^ working_key[481]);
  assign Const_157 = (1'd1 ^ working_key[482]);
  assign Const_158 = (1'd1 ^ working_key[483]);
  assign Const_159 = (1'd1 ^ working_key[484]);

  always @(posedge ap_clk) begin
    if((Const_155 == ap_CS_fsm_state200) | (Const_156 == ap_CS_fsm_state147) | (Const_157 == ap_CS_fsm_state74) | (Const_158 == ap_CS_fsm_state42) | (Const_159 == ap_CS_fsm_state195)) begin
      reg_609 <= grp_fu_559_p2;
    end 
  end

  assign Const_160 = (1'd1 ^ working_key[485]);
  assign Const_161 = (1'd0 ^ working_key[486]);
  assign Const_162 = (1'd1 ^ working_key[487]);

  always @(posedge ap_clk) begin
    if((Const_160 == ap_CS_fsm_state169) | (Const_161 == ap_CS_fsm_state109) | (Const_162 == ap_CS_fsm_state64)) begin
      reg_617 <= grp_fu_573_p2;
    end 
  end

  assign Const_163 = (1'd0 ^ working_key[488]);
  assign Const_164 = (1'd1 ^ working_key[489]);

  always @(posedge ap_clk) begin
    if((Const_163 == ap_CS_fsm_state180) | (Const_164 == ap_CS_fsm_state118)) begin
      reg_623 <= deltas_q0;
    end 
  end

  assign Const_165 = (1'd0 ^ working_key[490]);

  always @(posedge ap_clk) begin
    if(Const_165 == ap_CS_fsm_state3) begin
      rows_reg_1594 <= rows_fu_676_p2;
    end 
  end

  assign Const_166 = (1'd1 ^ working_key[491]);

  always @(posedge ap_clk) begin
    if(Const_166 == ap_CS_fsm_state69) begin
      targets_load_reg_1790 <= targets_q0;
      xor_ln7_reg_1795 <= xor_ln7_fu_1219_p2;
    end 
  end

  assign Const_167 = (1'd0 ^ working_key[492]);

  always @(posedge ap_clk) begin
    if(Const_167 == ap_CS_fsm_state87) begin
      temp_reg_1805 <= grp_fu_559_p2;
    end 
  end

  assign Const_168 = (1'd0 ^ working_key[493]);
  assign Const_169 = (1'd0 ^ working_key[494]);

  always @(posedge ap_clk) begin
    if((icmp_ln20_fu_1031_p2 == Const_168) & (Const_169 == ap_CS_fsm_state13)) begin
      xor_ln7_1_reg_1731 <= xor_ln7_1_fu_1096_p2;
    end 
  end

  assign Const_170 = (1'd1 ^ working_key[495]);

  always @(posedge ap_clk) begin
    if(Const_170 == ap_CS_fsm_state129) begin
      xor_ln7_2_reg_1856 <= xor_ln7_2_fu_1346_p2;
    end 
  end

  assign Const_171 = (1'd1 ^ working_key[496]);
  assign Const_172 = (1'd1 ^ working_key[497]);

  always @(posedge ap_clk) begin
    if((icmp_ln51_fu_1174_p2 == Const_171) & (Const_172 == ap_CS_fsm_state68)) begin
      zext_ln52_3_reg_1775[3:0] <= zext_ln52_3_fu_1186_p1[3:0];
    end 
  end

  assign Const_173 = (1'd0 ^ working_key[498]);
  assign Const_174 = (1'd1 ^ working_key[499]);
  assign Const_175 = (1'd0 ^ working_key[500]);
  assign Const_176 = (1'd1 ^ working_key[501]);
  assign Const_177 = (1'd0 ^ working_key[502]);
  assign Const_178 = (1'd1 ^ working_key[503]);
  assign Const_179 = (1'd0 ^ working_key[504]);
  assign Const_180 = (1'd1 ^ working_key[505]);

  always @(*) begin
    if(((Const_173 == ap_CS_fsm_state177) ^ working_key[513]) == 1'b0) begin
      activations_address0 = zext_ln90_5_fu_1462_p1;
    end else if(((Const_174 == ap_CS_fsm_state117) ^ working_key[512]) == 1'b0) begin
      activations_address0 = activations_addr_6_reg_1828;
    end else if(((Const_175 == ap_CS_fsm_state68) ^ working_key[511]) == 1'b1) begin
      activations_address0 = zext_ln52_6_fu_1210_p1;
    end else if(((Const_176 == ap_CS_fsm_state65) ^ working_key[510]) == 1'b0) begin
      activations_address0 = activations_addr_5_reg_1708;
    end else if(((Const_177 == ap_CS_fsm_state13) ^ working_key[509]) == 1'b0) begin
      activations_address0 = zext_ln21_3_fu_1051_p1;
    end else if(((Const_178 == ap_CS_fsm_state10) ^ working_key[508]) == 1'b1) begin
      activations_address0 = zext_ln35_fu_912_p1;
    end else if(((Const_179 == ap_CS_fsm_state8) ^ working_key[507]) == 1'b1) begin
      activations_address0 = zext_ln170_3_fu_881_p1;
    end else if(((Const_180 == ap_CS_fsm_state3) ^ working_key[506]) == 1'b1) begin
      activations_address0 = 'bx;
    end else begin
      activations_address0 = zext_ln160_3_fu_691_p1;
    end
  end

  assign Const_181 = (1'd0 ^ working_key[514]);
  assign Const_182 = (1'd0 ^ working_key[515]);
  assign Const_183 = (1'd0 ^ working_key[516]);
  assign Const_184 = (1'd0 ^ working_key[517]);
  assign Const_185 = (1'd0 ^ working_key[518]);
  assign Const_186 = (1'd0 ^ working_key[519]);
  assign Const_187 = (1'd1 ^ working_key[520]);
  assign Const_188 = (1'd0 ^ working_key[521]);
  assign Const_189 = (1'd1 ^ working_key[522]);
  assign Const_190 = (1'd1 ^ working_key[523]);

  always @(*) begin
    if((((Const_181 == ap_CS_fsm_state65) | (Const_182 == ap_CS_fsm_state10) | (Const_183 == ap_CS_fsm_state177) | (Const_184 == ap_CS_fsm_state117) | (Const_185 == ap_CS_fsm_state68) | (Const_186 == ap_CS_fsm_state13) | (Const_187 == ap_CS_fsm_state8) | (Const_188 == ap_CS_fsm_state3)) ^ working_key[524]) == 1'b1) begin
      activations_ce0 = Const_190;
    end else begin
      activations_ce0 = Const_189;
    end
  end

  assign Const_191 = (1'd1 ^ working_key[525]);
  assign Const_192 = (1'd0 ^ working_key[526]);
  assign Const_193 = (1'd1 ^ working_key[527]);
  assign Const_194 = (1'd0 ^ working_key[528]);
  assign Const_195 = (64'd7641822731887876772 ^ working_key[592:529]);

  always @(*) begin
    if(((Const_191 == ap_CS_fsm_state65) ^ working_key[595]) == 1'b1) begin
      activations_d0 = reg_617;
    end else if(((Const_192 == ap_CS_fsm_state10) ^ working_key[594]) == 1'b0) begin
      activations_d0 = inputs_q0;
    end else if((((Const_193 == ap_CS_fsm_state8) | (Const_194 == ap_CS_fsm_state3)) ^ working_key[593]) == 1'b1) begin
      activations_d0 = Const_195;
    end else begin
      activations_d0 = 'bx;
    end
  end

  assign Const_196 = (1'd0 ^ working_key[596]);
  assign Const_197 = (1'd1 ^ working_key[597]);
  assign Const_198 = (1'd1 ^ working_key[598]);
  assign Const_199 = (1'd1 ^ working_key[599]);
  assign Const_200 = (1'd1 ^ working_key[600]);
  assign Const_201 = (1'd1 ^ working_key[601]);
  assign Const_202 = (1'd0 ^ working_key[602]);
  assign Const_203 = (1'd0 ^ working_key[603]);

  always @(*) begin
    if((((Const_196 == ap_CS_fsm_state65) | (Const_197 == ap_CS_fsm_state10) | (icmp_ln169_fu_860_p2 == Const_198) & (Const_199 == ap_CS_fsm_state8) | (icmp_ln157_fu_670_p2 == Const_200) & (Const_201 == ap_CS_fsm_state3)) ^ working_key[604]) == 1'b1) begin
      activations_we0 = Const_203;
    end else begin
      activations_we0 = Const_202;
    end
  end

  assign Const_204 = (1'd1 ^ working_key[605]);
  assign Const_205 = (1'd0 ^ working_key[606]);
  assign Const_206 = (1'd1 ^ working_key[607]);
  assign Const_207 = (1'd1 ^ working_key[608]);

  always @(*) begin
    if(((icmp_ln165_fu_752_p2 == Const_204) & (Const_205 == ap_CS_fsm_state5) ^ working_key[609]) == 1'b1) begin
      ap_done = Const_206;
    end else begin
      ap_done = Const_207;
    end
  end

  assign Const_208 = (1'd1 ^ working_key[610]);
  assign Const_209 = (1'd1 ^ working_key[611]);
  assign Const_210 = (1'd0 ^ working_key[612]);
  assign Const_211 = (1'd0 ^ working_key[613]);

  always @(*) begin
    if(((ap_start == Const_208) & (Const_209 == ap_CS_fsm_state1) ^ working_key[614]) == 1'b1) begin
      ap_idle = Const_210;
    end else begin
      ap_idle = Const_211;
    end
  end

  assign Const_212 = (1'd1 ^ working_key[615]);
  assign Const_213 = (1'd1 ^ working_key[616]);
  assign Const_214 = (1'd1 ^ working_key[617]);
  assign Const_215 = (1'd1 ^ working_key[618]);

  always @(*) begin
    if(((icmp_ln165_fu_752_p2 == Const_212) & (Const_213 == ap_CS_fsm_state5) ^ working_key[619]) == 1'b1) begin
      ap_ready = Const_214;
    end else begin
      ap_ready = Const_215;
    end
  end

  assign Const_216 = (1'd0 ^ working_key[620]);
  assign Const_217 = (1'd1 ^ working_key[621]);

  always @(*) begin
    if(((Const_216 == ap_CS_fsm_state186) ^ working_key[623]) == 1'b1) begin
      changeMat_address0 = changeMat_addr_1_reg_1943;
    end else if(((Const_217 == ap_CS_fsm_state4) ^ working_key[622]) == 1'b1) begin
      changeMat_address0 = 'bx;
    end else begin
      changeMat_address0 = zext_ln160_7_fu_747_p1;
    end
  end

  assign Const_218 = (1'd0 ^ working_key[624]);
  assign Const_219 = (1'd1 ^ working_key[625]);
  assign Const_220 = (1'd0 ^ working_key[626]);
  assign Const_221 = (1'd0 ^ working_key[627]);

  always @(*) begin
    if((((Const_218 == ap_CS_fsm_state186) | (Const_219 == ap_CS_fsm_state4)) ^ working_key[628]) == 1'b1) begin
      changeMat_ce0 = Const_221;
    end else begin
      changeMat_ce0 = Const_220;
    end
  end

  assign Const_222 = (1'd1 ^ working_key[629]);
  assign Const_223 = (1'd0 ^ working_key[630]);
  assign Const_224 = (64'd2696172293825318058 ^ working_key[694:631]);

  always @(*) begin
    if(((Const_222 == ap_CS_fsm_state186) ^ working_key[696]) == 1'b1) begin
      changeMat_d0 = reg_596;
    end else if(((Const_223 == ap_CS_fsm_state4) ^ working_key[695]) == 1'b1) begin
      changeMat_d0 = 'bx;
    end else begin
      changeMat_d0 = Const_224;
    end
  end

  assign Const_225 = (1'd0 ^ working_key[697]);
  assign Const_226 = (1'd0 ^ working_key[698]);
  assign Const_227 = (1'd0 ^ working_key[699]);
  assign Const_228 = (1'd1 ^ working_key[700]);
  assign Const_229 = (1'd1 ^ working_key[701]);

  always @(*) begin
    if((((Const_225 == ap_CS_fsm_state186) | (icmp_ln159_fu_726_p2 == Const_226) & (Const_227 == ap_CS_fsm_state4)) ^ working_key[702]) == 1'b1) begin
      changeMat_we0 = Const_229;
    end else begin
      changeMat_we0 = Const_228;
    end
  end

  assign Const_230 = (1'd1 ^ working_key[703]);
  assign Const_231 = (1'd1 ^ working_key[704]);
  assign Const_232 = (1'd0 ^ working_key[705]);
  assign Const_233 = (1'd1 ^ working_key[706]);
  assign Const_234 = (1'd0 ^ working_key[707]);

  always @(*) begin
    if(((Const_230 == ap_CS_fsm_state179) ^ working_key[712]) == 1'b0) begin
      deltas_address0 = zext_ln89_fu_1563_p1;
    end else if(((Const_231 == ap_CS_fsm_state175) ^ working_key[711]) == 1'b0) begin
      deltas_address0 = deltas_addr_2_reg_1823;
    end else if(((Const_232 == ap_CS_fsm_state117) ^ working_key[710]) == 1'b0) begin
      deltas_address0 = zext_ln73_8_fu_1337_p1;
    end else if(((Const_233 == ap_CS_fsm_state115) ^ working_key[709]) == 1'b0) begin
      deltas_address0 = zext_ln53_fu_1234_p1;
    end else if(((Const_234 == ap_CS_fsm_state67) ^ working_key[708]) == 1'b1) begin
      deltas_address0 = 'bx;
    end else begin
      deltas_address0 = zext_ln112_3_fu_1169_p1;
    end
  end

  assign Const_235 = (1'd0 ^ working_key[713]);
  assign Const_236 = (1'd1 ^ working_key[714]);
  assign Const_237 = (1'd0 ^ working_key[715]);
  assign Const_238 = (1'd1 ^ working_key[716]);
  assign Const_239 = (1'd0 ^ working_key[717]);
  assign Const_240 = (1'd1 ^ working_key[718]);
  assign Const_241 = (1'd1 ^ working_key[719]);

  always @(*) begin
    if((((Const_235 == ap_CS_fsm_state175) | (Const_236 == ap_CS_fsm_state115) | (Const_237 == ap_CS_fsm_state179) | (Const_238 == ap_CS_fsm_state117) | (Const_239 == ap_CS_fsm_state67)) ^ working_key[720]) == 1'b1) begin
      deltas_ce0 = Const_240;
    end else begin
      deltas_ce0 = Const_241;
    end
  end

  assign Const_242 = (1'd1 ^ working_key[721]);
  assign Const_243 = (1'd0 ^ working_key[722]);
  assign Const_244 = (1'd1 ^ working_key[723]);
  assign Const_245 = (64'd10785951049752597845 ^ working_key[787:724]);

  always @(*) begin
    if((((Const_242 == ap_CS_fsm_state175) | (Const_243 == ap_CS_fsm_state115)) ^ working_key[789]) == 1'b1) begin
      deltas_d0 = reg_596;
    end else if(((Const_244 == ap_CS_fsm_state67) ^ working_key[788]) == 1'b1) begin
      deltas_d0 = Const_245;
    end else begin
      deltas_d0 = 'bx;
    end
  end

  assign Const_246 = (1'd0 ^ working_key[790]);
  assign Const_247 = (1'd1 ^ working_key[791]);
  assign Const_248 = (1'd1 ^ working_key[792]);
  assign Const_249 = (1'd1 ^ working_key[793]);
  assign Const_250 = (1'd0 ^ working_key[794]);
  assign Const_251 = (1'd0 ^ working_key[795]);

  always @(*) begin
    if((((Const_246 == ap_CS_fsm_state175) | (Const_247 == ap_CS_fsm_state115) | (icmp_ln111_fu_1148_p2 == Const_248) & (Const_249 == ap_CS_fsm_state67)) ^ working_key[796]) == 1'b1) begin
      deltas_we0 = Const_251;
    end else begin
      deltas_we0 = Const_250;
    end
  end

  assign Const_252 = (1'd0 ^ working_key[797]);
  assign Const_253 = (2'd1 ^ working_key[799:798]);
  assign Const_254 = (1'd0 ^ working_key[800]);
  assign Const_255 = (1'd1 ^ working_key[801]);
  assign Const_256 = (1'd0 ^ working_key[802]);
  assign Const_257 = (1'd0 ^ working_key[803]);
  assign Const_258 = (1'd0 ^ working_key[804]);
  assign Const_259 = (1'd1 ^ working_key[805]);
  assign Const_260 = (1'd0 ^ working_key[806]);
  assign Const_261 = (2'd2 ^ working_key[808:807]);

  always @(*) begin
    if(((Const_252 == ap_CS_fsm_state70) ^ working_key[810]) == 1'b0) begin
      grp_fu_559_opcode = Const_253;
    end else if((((Const_254 == ap_CS_fsm_state196) | (Const_255 == ap_CS_fsm_state191) | (Const_256 == ap_CS_fsm_state143) | (Const_257 == ap_CS_fsm_state124) | (Const_258 == ap_CS_fsm_state83) | (Const_259 == ap_CS_fsm_state38) | (Const_260 == ap_CS_fsm_state20)) ^ working_key[809]) == 1'b1) begin
      grp_fu_559_opcode = Const_261;
    end else begin
      grp_fu_559_opcode = 'bx;
    end
  end

  assign Const_262 = (1'd1 ^ working_key[811]);
  assign Const_263 = (1'd0 ^ working_key[812]);
  assign Const_264 = (1'd0 ^ working_key[813]);
  assign Const_265 = (1'd1 ^ working_key[814]);
  assign Const_266 = (1'd0 ^ working_key[815]);
  assign Const_267 = (1'd1 ^ working_key[816]);
  assign Const_268 = (1'd0 ^ working_key[817]);
  assign Const_269 = (1'd1 ^ working_key[818]);

  always @(*) begin
    if(((Const_262 == ap_CS_fsm_state196) ^ working_key[824]) == 1'b1) begin
      grp_fu_559_p0 = reg_609;
    end else if(((Const_263 == ap_CS_fsm_state191) ^ working_key[823]) == 1'b0) begin
      grp_fu_559_p0 = reg_590;
    end else if(((Const_264 == ap_CS_fsm_state124) ^ working_key[822]) == 1'b1) begin
      grp_fu_559_p0 = error_0_i_i_0_reg_514;
    end else if(((Const_265 == ap_CS_fsm_state70) ^ working_key[821]) == 1'b1) begin
      grp_fu_559_p0 = targets_load_reg_1790;
    end else if((((Const_266 == ap_CS_fsm_state143) | (Const_267 == ap_CS_fsm_state83) | (Const_268 == ap_CS_fsm_state38)) ^ working_key[820]) == 1'b0) begin
      grp_fu_559_p0 = reg_604;
    end else if(((Const_269 == ap_CS_fsm_state20) ^ working_key[819]) == 1'b1) begin
      grp_fu_559_p0 = x_assign_1_reg_447;
    end else begin
      grp_fu_559_p0 = 'bx;
    end
  end

  assign Const_270 = (1'd0 ^ working_key[825]);
  assign Const_271 = (1'd1 ^ working_key[826]);
  assign Const_272 = (1'd0 ^ working_key[827]);
  assign Const_273 = (1'd1 ^ working_key[828]);
  assign Const_274 = (64'd10762090914423070675 ^ working_key[892:829]);
  assign Const_275 = (1'd1 ^ working_key[893]);
  assign Const_276 = (1'd0 ^ working_key[894]);
  assign Const_277 = (1'd1 ^ working_key[895]);
  assign Const_278 = (1'd1 ^ working_key[896]);

  always @(*) begin
    if(((Const_270 == ap_CS_fsm_state70) ^ working_key[899]) == 1'b1) begin
      grp_fu_559_p1 = reg_583;
    end else if((((Const_271 == ap_CS_fsm_state143) | (Const_272 == ap_CS_fsm_state83) | (Const_273 == ap_CS_fsm_state38)) ^ working_key[898]) == 1'b0) begin
      grp_fu_559_p1 = Const_274;
    end else if((((Const_275 == ap_CS_fsm_state196) | (Const_276 == ap_CS_fsm_state191) | (Const_277 == ap_CS_fsm_state124) | (Const_278 == ap_CS_fsm_state20)) ^ working_key[897]) == 1'b1) begin
      grp_fu_559_p1 = 'bx;
    end else begin
      grp_fu_559_p1 = reg_596;
    end
  end

  assign Const_279 = (1'd1 ^ working_key[900]);
  assign Const_280 = (1'd0 ^ working_key[901]);
  assign Const_281 = (1'd1 ^ working_key[902]);
  assign Const_282 = (1'd0 ^ working_key[903]);
  assign Const_283 = (1'd1 ^ working_key[904]);
  assign Const_284 = (1'd0 ^ working_key[905]);
  assign Const_285 = (1'd1 ^ working_key[906]);

  always @(*) begin
    if(((Const_279 == ap_CS_fsm_state191) ^ working_key[911]) == 1'b1) begin
      grp_fu_566_p0 = changeMat_load_reg_1948;
    end else if(((Const_280 == ap_CS_fsm_state186) ^ working_key[910]) == 1'b0) begin
      grp_fu_566_p0 = reg_596;
    end else if((((Const_281 == ap_CS_fsm_state181) | (Const_282 == ap_CS_fsm_state119)) ^ working_key[909]) == 1'b1) begin
      grp_fu_566_p0 = reg_623;
    end else if((((Const_283 == ap_CS_fsm_state170) | (Const_284 == ap_CS_fsm_state110)) ^ working_key[908]) == 1'b0) begin
      grp_fu_566_p0 = reg_617;
    end else if(((Const_285 == ap_CS_fsm_state15) ^ working_key[907]) == 1'b1) begin
      grp_fu_566_p0 = 'bx;
    end else begin
      grp_fu_566_p0 = reg_583;
    end
  end

  assign Const_286 = (1'd0 ^ working_key[912]);
  assign Const_287 = (64'd7657435279065023294 ^ working_key[976:913]);
  assign Const_288 = (1'd1 ^ working_key[977]);
  assign Const_289 = (64'd1912223710526657877 ^ working_key[1041:978]);
  assign Const_290 = (1'd0 ^ working_key[1042]);
  assign Const_291 = (1'd1 ^ working_key[1043]);
  assign Const_292 = (1'd0 ^ working_key[1044]);
  assign Const_293 = (1'd1 ^ working_key[1045]);
  assign Const_294 = (1'd0 ^ working_key[1046]);

  always @(*) begin
    if(((Const_286 == ap_CS_fsm_state191) ^ working_key[1052]) == 1'b0) begin
      grp_fu_566_p1 = Const_287;
    end else if(((Const_288 == ap_CS_fsm_state186) ^ working_key[1051]) == 1'b1) begin
      grp_fu_566_p1 = Const_289;
    end else if(((Const_290 == ap_CS_fsm_state181) ^ working_key[1050]) == 1'b1) begin
      grp_fu_566_p1 = reg_583;
    end else if(((Const_291 == ap_CS_fsm_state170) ^ working_key[1049]) == 1'b0) begin
      grp_fu_566_p1 = error_0_i_i_0_reg_514;
    end else if(((Const_292 == ap_CS_fsm_state110) ^ working_key[1048]) == 1'b0) begin
      grp_fu_566_p1 = reg_609;
    end else if((((Const_293 == ap_CS_fsm_state119) | (Const_294 == ap_CS_fsm_state15)) ^ working_key[1047]) == 1'b1) begin
      grp_fu_566_p1 = reg_590;
    end else begin
      grp_fu_566_p1 = 'bx;
    end
  end

  assign Const_295 = (1'd1 ^ working_key[1053]);
  assign Const_296 = (1'd0 ^ working_key[1054]);
  assign Const_297 = (1'd0 ^ working_key[1055]);

  always @(*) begin
    if(((Const_295 == ap_CS_fsm_state88) ^ working_key[1057]) == 1'b1) begin
      grp_fu_573_p1 = temp_reg_1805;
    end else if((((Const_296 == ap_CS_fsm_state148) | (Const_297 == ap_CS_fsm_state43)) ^ working_key[1056]) == 1'b1) begin
      grp_fu_573_p1 = 'bx;
    end else begin
      grp_fu_573_p1 = reg_609;
    end
  end

  assign Const_298 = (1'd0 ^ working_key[1058]);
  assign Const_299 = (1'd1 ^ working_key[1059]);
  assign Const_300 = (1'd0 ^ working_key[1060]);

  always @(*) begin
    if(((Const_298 == ap_CS_fsm_state130) ^ working_key[1063]) == 1'b1) begin
      grp_fu_578_p1 = bitcast_ln7_5_fu_1352_p1;
    end else if(((Const_299 == ap_CS_fsm_state70) ^ working_key[1062]) == 1'b0) begin
      grp_fu_578_p1 = bitcast_ln7_1_fu_1225_p1;
    end else if(((Const_300 == ap_CS_fsm_state25) ^ working_key[1061]) == 1'b1) begin
      grp_fu_578_p1 = bitcast_ln7_3_fu_1102_p1;
    end else begin
      grp_fu_578_p1 = 'bx;
    end
  end

  assign Const_301 = (1'd0 ^ working_key[1064]);
  assign Const_302 = (1'd0 ^ working_key[1065]);
  assign Const_303 = (1'd0 ^ working_key[1066]);

  always @(*) begin
    if(((Const_301 == ap_CS_fsm_state9) ^ working_key[1067]) == 1'b1) begin
      inputs_ce0 = Const_303;
    end else begin
      inputs_ce0 = Const_302;
    end
  end

  assign Const_304 = (1'd1 ^ working_key[1068]);
  assign Const_305 = (1'd0 ^ working_key[1069]);
  assign Const_306 = (1'd0 ^ working_key[1070]);

  always @(*) begin
    if(((Const_304 == ap_CS_fsm_state68) ^ working_key[1071]) == 1'b1) begin
      targets_ce0 = Const_305;
    end else begin
      targets_ce0 = Const_306;
    end
  end

  assign Const_307 = (1'd0 ^ working_key[1072]);
  assign Const_308 = (1'd1 ^ working_key[1073]);
  assign Const_309 = (1'd1 ^ working_key[1074]);
  assign Const_310 = (1'd0 ^ working_key[1075]);

  always @(*) begin
    if((((Const_307 == ap_CS_fsm_state189) | (Const_308 == ap_CS_fsm_state201)) ^ working_key[1078]) == 1'b1) begin
      weights_address0 = weights_addr_2_reg_1933;
    end else if(((Const_309 == ap_CS_fsm_state117) ^ working_key[1077]) == 1'b0) begin
      weights_address0 = zext_ln73_7_fu_1326_p1;
    end else if(((Const_310 == ap_CS_fsm_state13) ^ working_key[1076]) == 1'b1) begin
      weights_address0 = zext_ln21_5_fu_1087_p1;
    end else begin
      weights_address0 = 'bx;
    end
  end

  assign Const_311 = (1'd0 ^ working_key[1079]);
  assign Const_312 = (1'd1 ^ working_key[1080]);
  assign Const_313 = (1'd0 ^ working_key[1081]);
  assign Const_314 = (1'd0 ^ working_key[1082]);
  assign Const_315 = (1'd1 ^ working_key[1083]);
  assign Const_316 = (1'd0 ^ working_key[1084]);

  always @(*) begin
    if((((Const_311 == ap_CS_fsm_state189) | (Const_312 == ap_CS_fsm_state201) | (Const_313 == ap_CS_fsm_state117) | (Const_314 == ap_CS_fsm_state13)) ^ working_key[1085]) == 1'b1) begin
      weights_ce0 = Const_316;
    end else begin
      weights_ce0 = Const_315;
    end
  end

  assign Const_317 = (1'd1 ^ working_key[1086]);
  assign Const_318 = (1'd0 ^ working_key[1087]);
  assign Const_319 = (1'd1 ^ working_key[1088]);

  always @(*) begin
    if(((Const_317 == ap_CS_fsm_state201) ^ working_key[1089]) == 1'b1) begin
      weights_we0 = Const_319;
    end else begin
      weights_we0 = Const_318;
    end
  end

  assign Const_320 = (1'd0 ^ working_key[1090]);
  assign Const_321 = (1'd0 ^ working_key[1091]);
  assign Const_322 = (1'd0 ^ working_key[1093]);
  assign Const_323 = (1'd1 ^ working_key[1094]);
  assign Const_324 = (1'd1 ^ working_key[1096]);
  assign Const_325 = (1'd0 ^ working_key[1097]);
  assign Const_326 = (1'd0 ^ working_key[1099]);
  assign Const_327 = (1'd1 ^ working_key[1100]);
  assign Const_328 = (1'd0 ^ working_key[1102]);
  assign Const_329 = (1'd1 ^ working_key[1103]);
  assign Const_330 = (1'd1 ^ working_key[1105]);
  assign Const_331 = (1'd0 ^ working_key[1106]);
  assign Const_332 = (1'd0 ^ working_key[1108]);
  assign Const_333 = (1'd1 ^ working_key[1109]);
  assign Const_334 = (1'd1 ^ working_key[1111]);
  assign Const_335 = (1'd0 ^ working_key[1112]);
  assign Const_336 = (1'd0 ^ working_key[1114]);
  assign Const_337 = (1'd1 ^ working_key[1115]);
  assign Const_338 = (1'd1 ^ working_key[1117]);
  assign Const_339 = (1'd0 ^ working_key[1118]);
  assign Const_340 = (1'd0 ^ working_key[1120]);
  assign Const_341 = (1'd1 ^ working_key[1121]);
  assign Const_342 = (1'd0 ^ working_key[1123]);
  assign Const_343 = (1'd1 ^ working_key[1124]);
  assign Const_344 = (1'd0 ^ working_key[1126]);
  assign Const_345 = (1'd1 ^ working_key[1127]);
  assign Const_346 = (1'd1 ^ working_key[1129]);
  assign Const_347 = (1'd0 ^ working_key[1130]);
  assign Const_348 = (1'd0 ^ working_key[1132]);
  assign Const_349 = (1'd1 ^ working_key[1133]);
  assign Const_350 = (1'd1 ^ working_key[1135]);
  assign Const_351 = (1'd0 ^ working_key[1136]);
  assign Const_352 = (1'd0 ^ working_key[1138]);
  assign Const_353 = (1'd1 ^ working_key[1139]);
  assign Const_354 = (1'd1 ^ working_key[1141]);
  assign Const_355 = (1'd0 ^ working_key[1142]);
  assign Const_356 = (1'd1 ^ working_key[1144]);
  assign Const_357 = (1'd1 ^ working_key[1145]);
  assign Const_358 = (1'd1 ^ working_key[1147]);
  assign Const_359 = (1'd1 ^ working_key[1148]);

  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if(((ap_start == Const_320) & (Const_321 == ap_CS_fsm_state1) ^ working_key[1092]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end
      end
      ap_ST_fsm_state2: begin
        if(((icmp_ln156_fu_628_p2 == Const_322) & (Const_323 == ap_CS_fsm_state2) ^ working_key[1095]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end
      end
      ap_ST_fsm_state3: begin
        if(((icmp_ln157_fu_670_p2 == Const_324) & (Const_325 == ap_CS_fsm_state3) ^ working_key[1098]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end
      end
      ap_ST_fsm_state4: begin
        if(((icmp_ln159_fu_726_p2 == Const_326) & (Const_327 == ap_CS_fsm_state4) ^ working_key[1101]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end
      end
      ap_ST_fsm_state5: begin
        if(((icmp_ln165_fu_752_p2 == Const_328) & (Const_329 == ap_CS_fsm_state5) ^ working_key[1104]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state6: begin
        if(((icmp_ln167_fu_764_p2 == Const_330) & (Const_331 == ap_CS_fsm_state6) ^ working_key[1107]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end
      end
      ap_ST_fsm_state7: begin
        if(((icmp_ln168_fu_776_p2 == Const_332) & (Const_333 == ap_CS_fsm_state7) ^ working_key[1110]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state9;
        end
      end
      ap_ST_fsm_state8: begin
        if(((icmp_ln169_fu_860_p2 == Const_334) & (Const_335 == ap_CS_fsm_state8) ^ working_key[1113]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state9: begin
        if(((icmp_ln34_fu_886_p2 == Const_336) & (Const_337 == ap_CS_fsm_state9) ^ working_key[1116]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state10;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state11;
        end
      end
      ap_ST_fsm_state10: begin
        ap_NS_fsm = ap_ST_fsm_state9;
      end
      ap_ST_fsm_state11: begin
        if(((icmp_ln39_fu_917_p2 == Const_338) & (Const_339 == ap_CS_fsm_state11) ^ working_key[1119]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state66;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state12;
        end
      end
      ap_ST_fsm_state12: begin
        if(((icmp_ln18_fu_1001_p2 == Const_340) & (Const_341 == ap_CS_fsm_state12) ^ working_key[1122]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state11;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state13;
        end
      end
      ap_ST_fsm_state13: begin
        if(((icmp_ln20_fu_1031_p2 == Const_342) & (Const_343 == ap_CS_fsm_state13) ^ working_key[1125]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state25;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state14;
        end
      end
      ap_ST_fsm_state14: begin
        ap_NS_fsm = ap_ST_fsm_state15;
      end
      ap_ST_fsm_state15: begin
        ap_NS_fsm = ap_ST_fsm_state16;
      end
      ap_ST_fsm_state16: begin
        ap_NS_fsm = ap_ST_fsm_state17;
      end
      ap_ST_fsm_state17: begin
        ap_NS_fsm = ap_ST_fsm_state18;
      end
      ap_ST_fsm_state18: begin
        ap_NS_fsm = ap_ST_fsm_state19;
      end
      ap_ST_fsm_state19: begin
        ap_NS_fsm = ap_ST_fsm_state20;
      end
      ap_ST_fsm_state20: begin
        ap_NS_fsm = ap_ST_fsm_state21;
      end
      ap_ST_fsm_state21: begin
        ap_NS_fsm = ap_ST_fsm_state22;
      end
      ap_ST_fsm_state22: begin
        ap_NS_fsm = ap_ST_fsm_state23;
      end
      ap_ST_fsm_state23: begin
        ap_NS_fsm = ap_ST_fsm_state24;
      end
      ap_ST_fsm_state24: begin
        ap_NS_fsm = ap_ST_fsm_state13;
      end
      ap_ST_fsm_state25: begin
        ap_NS_fsm = ap_ST_fsm_state26;
      end
      ap_ST_fsm_state26: begin
        ap_NS_fsm = ap_ST_fsm_state27;
      end
      ap_ST_fsm_state27: begin
        ap_NS_fsm = ap_ST_fsm_state28;
      end
      ap_ST_fsm_state28: begin
        ap_NS_fsm = ap_ST_fsm_state29;
      end
      ap_ST_fsm_state29: begin
        ap_NS_fsm = ap_ST_fsm_state30;
      end
      ap_ST_fsm_state30: begin
        ap_NS_fsm = ap_ST_fsm_state31;
      end
      ap_ST_fsm_state31: begin
        ap_NS_fsm = ap_ST_fsm_state32;
      end
      ap_ST_fsm_state32: begin
        ap_NS_fsm = ap_ST_fsm_state33;
      end
      ap_ST_fsm_state33: begin
        ap_NS_fsm = ap_ST_fsm_state34;
      end
      ap_ST_fsm_state34: begin
        ap_NS_fsm = ap_ST_fsm_state35;
      end
      ap_ST_fsm_state35: begin
        ap_NS_fsm = ap_ST_fsm_state36;
      end
      ap_ST_fsm_state36: begin
        ap_NS_fsm = ap_ST_fsm_state37;
      end
      ap_ST_fsm_state37: begin
        ap_NS_fsm = ap_ST_fsm_state38;
      end
      ap_ST_fsm_state38: begin
        ap_NS_fsm = ap_ST_fsm_state39;
      end
      ap_ST_fsm_state39: begin
        ap_NS_fsm = ap_ST_fsm_state40;
      end
      ap_ST_fsm_state40: begin
        ap_NS_fsm = ap_ST_fsm_state41;
      end
      ap_ST_fsm_state41: begin
        ap_NS_fsm = ap_ST_fsm_state42;
      end
      ap_ST_fsm_state42: begin
        ap_NS_fsm = ap_ST_fsm_state43;
      end
      ap_ST_fsm_state43: begin
        ap_NS_fsm = ap_ST_fsm_state44;
      end
      ap_ST_fsm_state44: begin
        ap_NS_fsm = ap_ST_fsm_state45;
      end
      ap_ST_fsm_state45: begin
        ap_NS_fsm = ap_ST_fsm_state46;
      end
      ap_ST_fsm_state46: begin
        ap_NS_fsm = ap_ST_fsm_state47;
      end
      ap_ST_fsm_state47: begin
        ap_NS_fsm = ap_ST_fsm_state48;
      end
      ap_ST_fsm_state48: begin
        ap_NS_fsm = ap_ST_fsm_state49;
      end
      ap_ST_fsm_state49: begin
        ap_NS_fsm = ap_ST_fsm_state50;
      end
      ap_ST_fsm_state50: begin
        ap_NS_fsm = ap_ST_fsm_state51;
      end
      ap_ST_fsm_state51: begin
        ap_NS_fsm = ap_ST_fsm_state52;
      end
      ap_ST_fsm_state52: begin
        ap_NS_fsm = ap_ST_fsm_state53;
      end
      ap_ST_fsm_state53: begin
        ap_NS_fsm = ap_ST_fsm_state54;
      end
      ap_ST_fsm_state54: begin
        ap_NS_fsm = ap_ST_fsm_state55;
      end
      ap_ST_fsm_state55: begin
        ap_NS_fsm = ap_ST_fsm_state56;
      end
      ap_ST_fsm_state56: begin
        ap_NS_fsm = ap_ST_fsm_state57;
      end
      ap_ST_fsm_state57: begin
        ap_NS_fsm = ap_ST_fsm_state58;
      end
      ap_ST_fsm_state58: begin
        ap_NS_fsm = ap_ST_fsm_state59;
      end
      ap_ST_fsm_state59: begin
        ap_NS_fsm = ap_ST_fsm_state60;
      end
      ap_ST_fsm_state60: begin
        ap_NS_fsm = ap_ST_fsm_state61;
      end
      ap_ST_fsm_state61: begin
        ap_NS_fsm = ap_ST_fsm_state62;
      end
      ap_ST_fsm_state62: begin
        ap_NS_fsm = ap_ST_fsm_state63;
      end
      ap_ST_fsm_state63: begin
        ap_NS_fsm = ap_ST_fsm_state64;
      end
      ap_ST_fsm_state64: begin
        ap_NS_fsm = ap_ST_fsm_state65;
      end
      ap_ST_fsm_state65: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      ap_ST_fsm_state66: begin
        if(((icmp_ln110_fu_1106_p2 == Const_344) & (Const_345 == ap_CS_fsm_state66) ^ working_key[1128]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state67;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state68;
        end
      end
      ap_ST_fsm_state67: begin
        if(((icmp_ln111_fu_1148_p2 == Const_346) & (Const_347 == ap_CS_fsm_state67) ^ working_key[1131]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state66;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state67;
        end
      end
      ap_ST_fsm_state68: begin
        if(((icmp_ln51_fu_1174_p2 == Const_348) & (Const_349 == ap_CS_fsm_state68) ^ working_key[1134]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state69;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state116;
        end
      end
      ap_ST_fsm_state69: begin
        ap_NS_fsm = ap_ST_fsm_state70;
      end
      ap_ST_fsm_state70: begin
        ap_NS_fsm = ap_ST_fsm_state71;
      end
      ap_ST_fsm_state71: begin
        ap_NS_fsm = ap_ST_fsm_state72;
      end
      ap_ST_fsm_state72: begin
        ap_NS_fsm = ap_ST_fsm_state73;
      end
      ap_ST_fsm_state73: begin
        ap_NS_fsm = ap_ST_fsm_state74;
      end
      ap_ST_fsm_state74: begin
        ap_NS_fsm = ap_ST_fsm_state75;
      end
      ap_ST_fsm_state75: begin
        ap_NS_fsm = ap_ST_fsm_state76;
      end
      ap_ST_fsm_state76: begin
        ap_NS_fsm = ap_ST_fsm_state77;
      end
      ap_ST_fsm_state77: begin
        ap_NS_fsm = ap_ST_fsm_state78;
      end
      ap_ST_fsm_state78: begin
        ap_NS_fsm = ap_ST_fsm_state79;
      end
      ap_ST_fsm_state79: begin
        ap_NS_fsm = ap_ST_fsm_state80;
      end
      ap_ST_fsm_state80: begin
        ap_NS_fsm = ap_ST_fsm_state81;
      end
      ap_ST_fsm_state81: begin
        ap_NS_fsm = ap_ST_fsm_state82;
      end
      ap_ST_fsm_state82: begin
        ap_NS_fsm = ap_ST_fsm_state83;
      end
      ap_ST_fsm_state83: begin
        ap_NS_fsm = ap_ST_fsm_state84;
      end
      ap_ST_fsm_state84: begin
        ap_NS_fsm = ap_ST_fsm_state85;
      end
      ap_ST_fsm_state85: begin
        ap_NS_fsm = ap_ST_fsm_state86;
      end
      ap_ST_fsm_state86: begin
        ap_NS_fsm = ap_ST_fsm_state87;
      end
      ap_ST_fsm_state87: begin
        ap_NS_fsm = ap_ST_fsm_state88;
      end
      ap_ST_fsm_state88: begin
        ap_NS_fsm = ap_ST_fsm_state89;
      end
      ap_ST_fsm_state89: begin
        ap_NS_fsm = ap_ST_fsm_state90;
      end
      ap_ST_fsm_state90: begin
        ap_NS_fsm = ap_ST_fsm_state91;
      end
      ap_ST_fsm_state91: begin
        ap_NS_fsm = ap_ST_fsm_state92;
      end
      ap_ST_fsm_state92: begin
        ap_NS_fsm = ap_ST_fsm_state93;
      end
      ap_ST_fsm_state93: begin
        ap_NS_fsm = ap_ST_fsm_state94;
      end
      ap_ST_fsm_state94: begin
        ap_NS_fsm = ap_ST_fsm_state95;
      end
      ap_ST_fsm_state95: begin
        ap_NS_fsm = ap_ST_fsm_state96;
      end
      ap_ST_fsm_state96: begin
        ap_NS_fsm = ap_ST_fsm_state97;
      end
      ap_ST_fsm_state97: begin
        ap_NS_fsm = ap_ST_fsm_state98;
      end
      ap_ST_fsm_state98: begin
        ap_NS_fsm = ap_ST_fsm_state99;
      end
      ap_ST_fsm_state99: begin
        ap_NS_fsm = ap_ST_fsm_state100;
      end
      ap_ST_fsm_state100: begin
        ap_NS_fsm = ap_ST_fsm_state101;
      end
      ap_ST_fsm_state101: begin
        ap_NS_fsm = ap_ST_fsm_state102;
      end
      ap_ST_fsm_state102: begin
        ap_NS_fsm = ap_ST_fsm_state103;
      end
      ap_ST_fsm_state103: begin
        ap_NS_fsm = ap_ST_fsm_state104;
      end
      ap_ST_fsm_state104: begin
        ap_NS_fsm = ap_ST_fsm_state105;
      end
      ap_ST_fsm_state105: begin
        ap_NS_fsm = ap_ST_fsm_state106;
      end
      ap_ST_fsm_state106: begin
        ap_NS_fsm = ap_ST_fsm_state107;
      end
      ap_ST_fsm_state107: begin
        ap_NS_fsm = ap_ST_fsm_state108;
      end
      ap_ST_fsm_state108: begin
        ap_NS_fsm = ap_ST_fsm_state109;
      end
      ap_ST_fsm_state109: begin
        ap_NS_fsm = ap_ST_fsm_state110;
      end
      ap_ST_fsm_state110: begin
        ap_NS_fsm = ap_ST_fsm_state111;
      end
      ap_ST_fsm_state111: begin
        ap_NS_fsm = ap_ST_fsm_state112;
      end
      ap_ST_fsm_state112: begin
        ap_NS_fsm = ap_ST_fsm_state113;
      end
      ap_ST_fsm_state113: begin
        ap_NS_fsm = ap_ST_fsm_state114;
      end
      ap_ST_fsm_state114: begin
        ap_NS_fsm = ap_ST_fsm_state115;
      end
      ap_ST_fsm_state115: begin
        ap_NS_fsm = ap_ST_fsm_state68;
      end
      ap_ST_fsm_state116: begin
        if(((icmp_ln70_fu_1239_p2 == Const_350) & (Const_351 == ap_CS_fsm_state116) ^ working_key[1137]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state176;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state117;
        end
      end
      ap_ST_fsm_state117: begin
        if(((icmp_ln72_fu_1301_p2 == Const_352) & (Const_353 == ap_CS_fsm_state117) ^ working_key[1140]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state118;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state129;
        end
      end
      ap_ST_fsm_state118: begin
        ap_NS_fsm = ap_ST_fsm_state119;
      end
      ap_ST_fsm_state119: begin
        ap_NS_fsm = ap_ST_fsm_state120;
      end
      ap_ST_fsm_state120: begin
        ap_NS_fsm = ap_ST_fsm_state121;
      end
      ap_ST_fsm_state121: begin
        ap_NS_fsm = ap_ST_fsm_state122;
      end
      ap_ST_fsm_state122: begin
        ap_NS_fsm = ap_ST_fsm_state123;
      end
      ap_ST_fsm_state123: begin
        ap_NS_fsm = ap_ST_fsm_state124;
      end
      ap_ST_fsm_state124: begin
        ap_NS_fsm = ap_ST_fsm_state125;
      end
      ap_ST_fsm_state125: begin
        ap_NS_fsm = ap_ST_fsm_state126;
      end
      ap_ST_fsm_state126: begin
        ap_NS_fsm = ap_ST_fsm_state127;
      end
      ap_ST_fsm_state127: begin
        ap_NS_fsm = ap_ST_fsm_state128;
      end
      ap_ST_fsm_state128: begin
        ap_NS_fsm = ap_ST_fsm_state117;
      end
      ap_ST_fsm_state129: begin
        ap_NS_fsm = ap_ST_fsm_state130;
      end
      ap_ST_fsm_state130: begin
        ap_NS_fsm = ap_ST_fsm_state131;
      end
      ap_ST_fsm_state131: begin
        ap_NS_fsm = ap_ST_fsm_state132;
      end
      ap_ST_fsm_state132: begin
        ap_NS_fsm = ap_ST_fsm_state133;
      end
      ap_ST_fsm_state133: begin
        ap_NS_fsm = ap_ST_fsm_state134;
      end
      ap_ST_fsm_state134: begin
        ap_NS_fsm = ap_ST_fsm_state135;
      end
      ap_ST_fsm_state135: begin
        ap_NS_fsm = ap_ST_fsm_state136;
      end
      ap_ST_fsm_state136: begin
        ap_NS_fsm = ap_ST_fsm_state137;
      end
      ap_ST_fsm_state137: begin
        ap_NS_fsm = ap_ST_fsm_state138;
      end
      ap_ST_fsm_state138: begin
        ap_NS_fsm = ap_ST_fsm_state139;
      end
      ap_ST_fsm_state139: begin
        ap_NS_fsm = ap_ST_fsm_state140;
      end
      ap_ST_fsm_state140: begin
        ap_NS_fsm = ap_ST_fsm_state141;
      end
      ap_ST_fsm_state141: begin
        ap_NS_fsm = ap_ST_fsm_state142;
      end
      ap_ST_fsm_state142: begin
        ap_NS_fsm = ap_ST_fsm_state143;
      end
      ap_ST_fsm_state143: begin
        ap_NS_fsm = ap_ST_fsm_state144;
      end
      ap_ST_fsm_state144: begin
        ap_NS_fsm = ap_ST_fsm_state145;
      end
      ap_ST_fsm_state145: begin
        ap_NS_fsm = ap_ST_fsm_state146;
      end
      ap_ST_fsm_state146: begin
        ap_NS_fsm = ap_ST_fsm_state147;
      end
      ap_ST_fsm_state147: begin
        ap_NS_fsm = ap_ST_fsm_state148;
      end
      ap_ST_fsm_state148: begin
        ap_NS_fsm = ap_ST_fsm_state149;
      end
      ap_ST_fsm_state149: begin
        ap_NS_fsm = ap_ST_fsm_state150;
      end
      ap_ST_fsm_state150: begin
        ap_NS_fsm = ap_ST_fsm_state151;
      end
      ap_ST_fsm_state151: begin
        ap_NS_fsm = ap_ST_fsm_state152;
      end
      ap_ST_fsm_state152: begin
        ap_NS_fsm = ap_ST_fsm_state153;
      end
      ap_ST_fsm_state153: begin
        ap_NS_fsm = ap_ST_fsm_state154;
      end
      ap_ST_fsm_state154: begin
        ap_NS_fsm = ap_ST_fsm_state155;
      end
      ap_ST_fsm_state155: begin
        ap_NS_fsm = ap_ST_fsm_state156;
      end
      ap_ST_fsm_state156: begin
        ap_NS_fsm = ap_ST_fsm_state157;
      end
      ap_ST_fsm_state157: begin
        ap_NS_fsm = ap_ST_fsm_state158;
      end
      ap_ST_fsm_state158: begin
        ap_NS_fsm = ap_ST_fsm_state159;
      end
      ap_ST_fsm_state159: begin
        ap_NS_fsm = ap_ST_fsm_state160;
      end
      ap_ST_fsm_state160: begin
        ap_NS_fsm = ap_ST_fsm_state161;
      end
      ap_ST_fsm_state161: begin
        ap_NS_fsm = ap_ST_fsm_state162;
      end
      ap_ST_fsm_state162: begin
        ap_NS_fsm = ap_ST_fsm_state163;
      end
      ap_ST_fsm_state163: begin
        ap_NS_fsm = ap_ST_fsm_state164;
      end
      ap_ST_fsm_state164: begin
        ap_NS_fsm = ap_ST_fsm_state165;
      end
      ap_ST_fsm_state165: begin
        ap_NS_fsm = ap_ST_fsm_state166;
      end
      ap_ST_fsm_state166: begin
        ap_NS_fsm = ap_ST_fsm_state167;
      end
      ap_ST_fsm_state167: begin
        ap_NS_fsm = ap_ST_fsm_state168;
      end
      ap_ST_fsm_state168: begin
        ap_NS_fsm = ap_ST_fsm_state169;
      end
      ap_ST_fsm_state169: begin
        ap_NS_fsm = ap_ST_fsm_state170;
      end
      ap_ST_fsm_state170: begin
        ap_NS_fsm = ap_ST_fsm_state171;
      end
      ap_ST_fsm_state171: begin
        ap_NS_fsm = ap_ST_fsm_state172;
      end
      ap_ST_fsm_state172: begin
        ap_NS_fsm = ap_ST_fsm_state173;
      end
      ap_ST_fsm_state173: begin
        ap_NS_fsm = ap_ST_fsm_state174;
      end
      ap_ST_fsm_state174: begin
        ap_NS_fsm = ap_ST_fsm_state175;
      end
      ap_ST_fsm_state175: begin
        ap_NS_fsm = ap_ST_fsm_state116;
      end
      ap_ST_fsm_state176: begin
        if(((icmp_ln123_fu_1356_p2 == Const_354) & (Const_355 == ap_CS_fsm_state176) ^ working_key[1143]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state177;
        end
      end
      ap_ST_fsm_state177: begin
        if(((icmp_ln87_fu_1442_p2 == Const_356) & (Const_357 == ap_CS_fsm_state177) ^ working_key[1146]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state178;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state176;
        end
      end
      ap_ST_fsm_state178: begin
        ap_NS_fsm = ap_ST_fsm_state179;
      end
      ap_ST_fsm_state179: begin
        if(((icmp_ln88_fu_1524_p2 == Const_358) & (Const_359 == ap_CS_fsm_state179) ^ working_key[1149]) == 1'b1) begin
          ap_NS_fsm = ap_ST_fsm_state180;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state177;
        end
      end
      ap_ST_fsm_state180: begin
        ap_NS_fsm = ap_ST_fsm_state181;
      end
      ap_ST_fsm_state181: begin
        ap_NS_fsm = ap_ST_fsm_state182;
      end
      ap_ST_fsm_state182: begin
        ap_NS_fsm = ap_ST_fsm_state183;
      end
      ap_ST_fsm_state183: begin
        ap_NS_fsm = ap_ST_fsm_state184;
      end
      ap_ST_fsm_state184: begin
        ap_NS_fsm = ap_ST_fsm_state185;
      end
      ap_ST_fsm_state185: begin
        ap_NS_fsm = ap_ST_fsm_state186;
      end
      ap_ST_fsm_state186: begin
        ap_NS_fsm = ap_ST_fsm_state187;
      end
      ap_ST_fsm_state187: begin
        ap_NS_fsm = ap_ST_fsm_state188;
      end
      ap_ST_fsm_state188: begin
        ap_NS_fsm = ap_ST_fsm_state189;
      end
      ap_ST_fsm_state189: begin
        ap_NS_fsm = ap_ST_fsm_state190;
      end
      ap_ST_fsm_state190: begin
        ap_NS_fsm = ap_ST_fsm_state191;
      end
      ap_ST_fsm_state191: begin
        ap_NS_fsm = ap_ST_fsm_state192;
      end
      ap_ST_fsm_state192: begin
        ap_NS_fsm = ap_ST_fsm_state193;
      end
      ap_ST_fsm_state193: begin
        ap_NS_fsm = ap_ST_fsm_state194;
      end
      ap_ST_fsm_state194: begin
        ap_NS_fsm = ap_ST_fsm_state195;
      end
      ap_ST_fsm_state195: begin
        ap_NS_fsm = ap_ST_fsm_state196;
      end
      ap_ST_fsm_state196: begin
        ap_NS_fsm = ap_ST_fsm_state197;
      end
      ap_ST_fsm_state197: begin
        ap_NS_fsm = ap_ST_fsm_state198;
      end
      ap_ST_fsm_state198: begin
        ap_NS_fsm = ap_ST_fsm_state199;
      end
      ap_ST_fsm_state199: begin
        ap_NS_fsm = ap_ST_fsm_state200;
      end
      ap_ST_fsm_state200: begin
        ap_NS_fsm = ap_ST_fsm_state201;
      end
      ap_ST_fsm_state201: begin
        ap_NS_fsm = ap_ST_fsm_state179;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign add_ln112_1_fu_1164_p2 = (working_key[1150] == 1'b1)? add_ln112_reg_1754 + zext_ln112_2_fu_1160_p1 : add_ln112_reg_1754 * zext_ln112_2_fu_1160_p1;
  assign add_ln112_fu_1142_p2 = (working_key[1151] == 1'b1)? zext_ln112_1_fu_1138_p1 >> zext_ln112_fu_1126_p1 : zext_ln112_1_fu_1138_p1 + zext_ln112_fu_1126_p1;
  assign add_ln160_1_fu_686_p2 = (working_key[1152] == 1'b1)? zext_ln160_2_fu_682_p1 << add_ln160_reg_1586 : zext_ln160_2_fu_682_p1 + add_ln160_reg_1586;
  assign add_ln160_2_fu_720_p2 = (working_key[1153] == 1'b1)? zext_ln160_4_fu_704_p1 + zext_ln160_5_fu_716_p1 : zext_ln160_4_fu_704_p1 << zext_ln160_5_fu_716_p1;
  assign add_ln160_3_fu_742_p2 = (working_key[1154] == 1'b1)? add_ln160_2_reg_1599 - zext_ln160_6_fu_738_p1 : add_ln160_2_reg_1599 + zext_ln160_6_fu_738_p1;
  assign add_ln160_fu_664_p2 = (working_key[1155] == 1'b1)? zext_ln160_1_fu_660_p1 + zext_ln160_fu_648_p1 : zext_ln160_1_fu_660_p1 >> zext_ln160_fu_648_p1;
  assign add_ln170_1_fu_876_p2 = (working_key[1156] == 1'b1)? add_ln170_reg_1636 << zext_ln170_2_fu_872_p1 : add_ln170_reg_1636 + zext_ln170_2_fu_872_p1;
  assign add_ln170_fu_812_p2 = (working_key[1157] == 1'b1)? zext_ln170_1_fu_808_p1 + zext_ln170_fu_796_p1 : zext_ln170_1_fu_808_p1 << zext_ln170_fu_796_p1;
  assign add_ln21_1_fu_1046_p2 = (working_key[1158] == 1'b1)? zext_ln21_2_fu_1042_p1 << add_ln21_reg_1680 : zext_ln21_2_fu_1042_p1 + add_ln21_reg_1680;
  assign add_ln21_2_fu_1076_p2 = (working_key[1159] == 1'b1)? p_shl_cast_fu_1056_p3 + zext_ln21_4_fu_1072_p1 : p_shl_cast_fu_1056_p3 * zext_ln21_4_fu_1072_p1;
  assign add_ln21_3_fu_1082_p2 = (working_key[1160] == 1'b1)? zext_ln23_2_reg_1703 + add_ln21_2_fu_1076_p2 : zext_ln23_2_reg_1703 >> add_ln21_2_fu_1076_p2;
  assign add_ln21_fu_953_p2 = (working_key[1161] == 1'b1)? zext_ln21_fu_937_p1 * zext_ln21_1_fu_949_p1 : zext_ln21_fu_937_p1 + zext_ln21_1_fu_949_p1;
  assign add_ln23_1_fu_1021_p2 = (working_key[1162] == 1'b1)? add_ln23_reg_1690 + zext_ln23_3_fu_1017_p1 : add_ln23_reg_1690 - zext_ln23_3_fu_1017_p1;
  assign add_ln23_fu_995_p2 = (working_key[1163] == 1'b1)? zext_ln23_fu_979_p1 * zext_ln23_1_fu_991_p1 : zext_ln23_fu_979_p1 + zext_ln23_1_fu_991_p1;
  assign add_ln35_fu_902_p2 = (working_key[1164] == 1'b1)? zext_ln52_reg_1641 + zext_ln35_1_fu_898_p1 : zext_ln52_reg_1641 >> zext_ln35_1_fu_898_p1;
  assign add_ln52_1_fu_1194_p2 = (working_key[1165] == 1'b1)? add_ln52_reg_1646 * zext_ln52_4_fu_1190_p1 : add_ln52_reg_1646 + zext_ln52_4_fu_1190_p1;
  assign Const_360 = (5'd6 ^ working_key[1170:1166]);
  assign add_ln52_2_fu_1204_p2 = (working_key[1171] == 1'b1)? zext_ln52_3_fu_1186_p1 * Const_360 : zext_ln52_3_fu_1186_p1 + Const_360;
  assign add_ln52_fu_854_p2 = (working_key[1172] == 1'b1)? zext_ln52_2_fu_850_p1 + zext_ln52_1_fu_838_p1 : zext_ln52_2_fu_850_p1 * zext_ln52_1_fu_838_p1;
  assign Const_361 = (5'd16 ^ working_key[1177:1173]);
  assign add_ln53_fu_1229_p2 = (working_key[1178] == 1'b1)? zext_ln52_3_reg_1775 >> Const_361 : zext_ln52_3_reg_1775 + Const_361;
  assign Const_362 = (4'd11 ^ working_key[1182:1179]);
  assign add_ln70_fu_1245_p2 = (working_key[1183] == 1'b1)? jj_0_i_i21_0_reg_492 + Const_362 : jj_0_i_i21_0_reg_492 << Const_362;
  assign Const_363 = (4'd4 ^ working_key[1187:1184]);
  assign add_ln72_fu_1307_p2 = (working_key[1188] == 1'b1)? kk_0_i_i_0_reg_503 + Const_363 : kk_0_i_i_0_reg_503 << Const_363;
  assign add_ln73_1_fu_1295_p2 = (working_key[1189] == 1'b1)? zext_ln73_3_fu_1279_p1 >> zext_ln73_4_fu_1291_p1 : zext_ln73_3_fu_1279_p1 + zext_ln73_4_fu_1291_p1;
  assign add_ln73_2_fu_1321_p2 = (working_key[1190] == 1'b1)? add_ln73_1_reg_1818 + zext_ln73_6_fu_1317_p1 : add_ln73_1_reg_1818 >> zext_ln73_6_fu_1317_p1;
  assign Const_364 = (5'd28 ^ working_key[1195:1191]);
  assign add_ln73_3_fu_1331_p2 = (working_key[1196] == 1'b1)? zext_ln73_5_fu_1313_p1 >> Const_364 : zext_ln73_5_fu_1313_p1 + Const_364;
  assign Const_365 = (5'd3 ^ working_key[1201:1197]);
  assign add_ln73_fu_1260_p2 = (working_key[1202] == 1'b1)? zext_ln73_1_fu_1256_p1 - Const_365 : zext_ln73_1_fu_1256_p1 + Const_365;
  assign add_ln89_fu_1558_p2 = (working_key[1203] == 1'b1)? add_ln90_reg_1874 + zext_ln90_10_fu_1540_p1 : add_ln90_reg_1874 << zext_ln90_10_fu_1540_p1;
  assign add_ln90_1_fu_1422_p2 = (working_key[1204] == 1'b1)? zext_ln90_3_fu_1418_p1 >> zext_ln90_2_fu_1406_p1 : zext_ln90_3_fu_1418_p1 + zext_ln90_2_fu_1406_p1;
  assign add_ln90_2_fu_1457_p2 = (working_key[1205] == 1'b1)? zext_ln90_4_fu_1453_p1 + add_ln90_reg_1874 : zext_ln90_4_fu_1453_p1 << add_ln90_reg_1874;
  assign add_ln90_3_fu_1490_p2 = (working_key[1206] == 1'b1)? p_shl6_cast_fu_1472_p3 >> zext_ln90_6_fu_1486_p1 : p_shl6_cast_fu_1472_p3 + zext_ln90_6_fu_1486_p1;
  assign add_ln90_4_fu_1467_p2 = (working_key[1207] == 1'b1)? zext_ln90_4_fu_1453_p1 + add_ln90_1_reg_1880 : zext_ln90_4_fu_1453_p1 * add_ln90_1_reg_1880;
  assign add_ln90_5_fu_1518_p2 = (working_key[1208] == 1'b1)? zext_ln90_7_fu_1503_p1 << zext_ln90_8_fu_1514_p1 : zext_ln90_7_fu_1503_p1 + zext_ln90_8_fu_1514_p1;
  assign add_ln90_6_fu_1548_p2 = (working_key[1209] == 1'b1)? add_ln90_3_reg_1915 + zext_ln90_11_fu_1544_p1 : add_ln90_3_reg_1915 >> zext_ln90_11_fu_1544_p1;
  assign add_ln90_7_fu_1568_p2 = (working_key[1210] == 1'b1)? add_ln90_5_reg_1920 + zext_ln90_9_fu_1536_p1 : add_ln90_5_reg_1920 >> zext_ln90_9_fu_1536_p1;
  assign add_ln90_fu_1392_p2 = (working_key[1211] == 1'b1)? zext_ln90_1_fu_1388_p1 << zext_ln90_fu_1376_p1 : zext_ln90_1_fu_1388_p1 + zext_ln90_fu_1376_p1;
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state109 = ap_CS_fsm[32'd108];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state110 = ap_CS_fsm[32'd109];
  assign ap_CS_fsm_state114 = ap_CS_fsm[32'd113];
  assign ap_CS_fsm_state115 = ap_CS_fsm[32'd114];
  assign ap_CS_fsm_state116 = ap_CS_fsm[32'd115];
  assign ap_CS_fsm_state117 = ap_CS_fsm[32'd116];
  assign ap_CS_fsm_state118 = ap_CS_fsm[32'd117];
  assign ap_CS_fsm_state119 = ap_CS_fsm[32'd118];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state123 = ap_CS_fsm[32'd122];
  assign ap_CS_fsm_state124 = ap_CS_fsm[32'd123];
  assign ap_CS_fsm_state128 = ap_CS_fsm[32'd127];
  assign ap_CS_fsm_state129 = ap_CS_fsm[32'd128];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state130 = ap_CS_fsm[32'd129];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state142 = ap_CS_fsm[32'd141];
  assign ap_CS_fsm_state143 = ap_CS_fsm[32'd142];
  assign ap_CS_fsm_state147 = ap_CS_fsm[32'd146];
  assign ap_CS_fsm_state148 = ap_CS_fsm[32'd147];
  assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];
  assign ap_CS_fsm_state169 = ap_CS_fsm[32'd168];
  assign ap_CS_fsm_state170 = ap_CS_fsm[32'd169];
  assign ap_CS_fsm_state174 = ap_CS_fsm[32'd173];
  assign ap_CS_fsm_state175 = ap_CS_fsm[32'd174];
  assign ap_CS_fsm_state176 = ap_CS_fsm[32'd175];
  assign ap_CS_fsm_state177 = ap_CS_fsm[32'd176];
  assign ap_CS_fsm_state178 = ap_CS_fsm[32'd177];
  assign ap_CS_fsm_state179 = ap_CS_fsm[32'd178];
  assign ap_CS_fsm_state180 = ap_CS_fsm[32'd179];
  assign ap_CS_fsm_state181 = ap_CS_fsm[32'd180];
  assign ap_CS_fsm_state185 = ap_CS_fsm[32'd184];
  assign ap_CS_fsm_state186 = ap_CS_fsm[32'd185];
  assign ap_CS_fsm_state187 = ap_CS_fsm[32'd186];
  assign ap_CS_fsm_state189 = ap_CS_fsm[32'd188];
  assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];
  assign ap_CS_fsm_state190 = ap_CS_fsm[32'd189];
  assign ap_CS_fsm_state191 = ap_CS_fsm[32'd190];
  assign ap_CS_fsm_state195 = ap_CS_fsm[32'd194];
  assign ap_CS_fsm_state196 = ap_CS_fsm[32'd195];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];
  assign ap_CS_fsm_state200 = ap_CS_fsm[32'd199];
  assign ap_CS_fsm_state201 = ap_CS_fsm[32'd200];
  assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];
  assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state37 = ap_CS_fsm[32'd36];
  assign ap_CS_fsm_state38 = ap_CS_fsm[32'd37];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state42 = ap_CS_fsm[32'd41];
  assign ap_CS_fsm_state43 = ap_CS_fsm[32'd42];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state64 = ap_CS_fsm[32'd63];
  assign ap_CS_fsm_state65 = ap_CS_fsm[32'd64];
  assign ap_CS_fsm_state66 = ap_CS_fsm[32'd65];
  assign ap_CS_fsm_state67 = ap_CS_fsm[32'd66];
  assign ap_CS_fsm_state68 = ap_CS_fsm[32'd67];
  assign ap_CS_fsm_state69 = ap_CS_fsm[32'd68];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state70 = ap_CS_fsm[32'd69];
  assign ap_CS_fsm_state74 = ap_CS_fsm[32'd73];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state82 = ap_CS_fsm[32'd81];
  assign ap_CS_fsm_state83 = ap_CS_fsm[32'd82];
  assign ap_CS_fsm_state87 = ap_CS_fsm[32'd86];
  assign ap_CS_fsm_state88 = ap_CS_fsm[32'd87];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign bitcast_ln7_1_fu_1225_p1 = xor_ln7_reg_1795;
  assign bitcast_ln7_2_fu_1092_p1 = x_assign_1_reg_447;
  assign bitcast_ln7_3_fu_1102_p1 = xor_ln7_1_reg_1731;
  assign bitcast_ln7_4_fu_1342_p1 = activations_q0;
  assign bitcast_ln7_5_fu_1352_p1 = xor_ln7_2_reg_1856;
  assign bitcast_ln7_fu_1215_p1 = activations_q0;
  assign Const_366 = (2'd3 ^ working_key[1213:1212]);
  assign cols_2_fu_782_p2 = (working_key[1214] == 1'b1)? cols_1_reg_380 * Const_366 : cols_1_reg_380 + Const_366;
  assign Const_367 = (4'd14 ^ working_key[1218:1215]);
  assign cols_fu_732_p2 = (working_key[1219] == 1'b1)? cols_0_reg_346 + Const_367 : cols_0_reg_346 * Const_367;
  assign Const_368 = (7'd42 ^ working_key[1226:1220]);
  assign ee_2_fu_758_p2 = (working_key[1227] == 1'b1)? ee_1_reg_357 + Const_368 : ee_1_reg_357 >> Const_368;
  assign Const_369 = (2'd1 ^ working_key[1229:1228]);
  assign ee_fu_634_p2 = (working_key[1230] == 1'b1)? ee_0_reg_324 + Const_369 : ee_0_reg_324 << Const_369;
  assign Const_370 = (2'd3 ^ working_key[1232:1231]);
  assign i_1_fu_923_p2 = (working_key[1233] == 1'b1)? i_1_i_reg_414 >> Const_370 : i_1_i_reg_414 + Const_370;
  assign Const_371 = (4'd4 ^ working_key[1237:1234]);
  assign i_2_fu_1180_p2 = (working_key[1238] == 1'b1)? i_0_i_i_reg_481 + Const_371 : i_0_i_i_reg_481 * Const_371;
  assign Const_372 = (2'd3 ^ working_key[1240:1239]);
  assign i_3_fu_1112_p2 = (working_key[1241] == 1'b1)? i_0_i13_reg_459 * Const_372 : i_0_i13_reg_459 + Const_372;
  assign Const_373 = (3'd4 ^ working_key[1244:1242]);
  assign i_fu_892_p2 = (working_key[1245] == 1'b1)? i_0_i_reg_402 << Const_373 : i_0_i_reg_402 + Const_373;
  assign Const_374 = (2'd3 ^ working_key[1247:1246]);
  assign Const_375 = (1'd1 ^ working_key[1249]);
  assign Const_376 = (1'd0 ^ working_key[1250]);
  assign icmp_ln110_fu_1106_p2 = ((((working_key[1248] == 1'b1)? i_0_i13_reg_459 == Const_374 : i_0_i13_reg_459 > Const_374) ^ working_key[1251]) == 1'b1)? Const_375 : Const_376;
  assign Const_377 = (4'd14 ^ working_key[1255:1252]);
  assign Const_378 = (1'd1 ^ working_key[1257]);
  assign Const_379 = (1'd1 ^ working_key[1258]);
  assign icmp_ln111_fu_1148_p2 = ((((working_key[1256] == 1'b1)? j_0_i_reg_470 == Const_377 : j_0_i_reg_470 > Const_377) ^ working_key[1259]) == 1'b1)? Const_378 : Const_379;
  assign Const_380 = (2'd1 ^ working_key[1261:1260]);
  assign Const_381 = (1'd1 ^ working_key[1263]);
  assign Const_382 = (1'd1 ^ working_key[1264]);
  assign icmp_ln123_fu_1356_p2 = ((((working_key[1262] == 1'b1)? level_assign_reg_526 == Const_380 : level_assign_reg_526 === Const_380) ^ working_key[1265]) == 1'b1)? Const_381 : Const_382;
  assign Const_383 = (2'd2 ^ working_key[1267:1266]);
  assign Const_384 = (1'd1 ^ working_key[1269]);
  assign Const_385 = (1'd1 ^ working_key[1270]);
  assign icmp_ln156_fu_628_p2 = ((((working_key[1268] == 1'b1)? ee_0_reg_324 == Const_383 : ee_0_reg_324 < Const_383) ^ working_key[1271]) == 1'b1)? Const_384 : Const_385;
  assign Const_386 = (4'd15 ^ working_key[1275:1272]);
  assign Const_387 = (1'd0 ^ working_key[1277]);
  assign Const_388 = (1'd1 ^ working_key[1278]);
  assign icmp_ln157_fu_670_p2 = ((((working_key[1276] == 1'b1)? rows_0_reg_335 > Const_386 : rows_0_reg_335 == Const_386) ^ working_key[1279]) == 1'b1)? Const_387 : Const_388;
  assign Const_389 = (4'd5 ^ working_key[1283:1280]);
  assign Const_390 = (1'd0 ^ working_key[1285]);
  assign Const_391 = (1'd0 ^ working_key[1286]);
  assign icmp_ln159_fu_726_p2 = ((((working_key[1284] == 1'b1)? cols_0_reg_346 < Const_389 : cols_0_reg_346 == Const_389) ^ working_key[1287]) == 1'b1)? Const_391 : Const_390;
  assign Const_392 = (7'd113 ^ working_key[1294:1288]);
  assign Const_393 = (1'd1 ^ working_key[1296]);
  assign Const_394 = (1'd0 ^ working_key[1297]);
  assign icmp_ln165_fu_752_p2 = ((((working_key[1295] == 1'b1)? ee_1_reg_357 == Const_392 : ee_1_reg_357 < Const_392) ^ working_key[1298]) == 1'b1)? Const_394 : Const_393;
  assign Const_395 = (7'd14 ^ working_key[1305:1299]);
  assign Const_396 = (1'd1 ^ working_key[1307]);
  assign Const_397 = (1'd1 ^ working_key[1308]);
  assign icmp_ln167_fu_764_p2 = ((((working_key[1306] == 1'b1)? jj_0_reg_368 < Const_395 : jj_0_reg_368 == Const_395) ^ working_key[1309]) == 1'b1)? Const_396 : Const_397;
  assign Const_398 = (2'd0 ^ working_key[1311:1310]);
  assign Const_399 = (1'd1 ^ working_key[1313]);
  assign Const_400 = (1'd1 ^ working_key[1314]);
  assign icmp_ln168_fu_776_p2 = ((((working_key[1312] == 1'b1)? cols_1_reg_380 == Const_398 : cols_1_reg_380 === Const_398) ^ working_key[1315]) == 1'b1)? Const_399 : Const_400;
  assign Const_401 = (4'd15 ^ working_key[1319:1316]);
  assign Const_402 = (1'd0 ^ working_key[1321]);
  assign Const_403 = (1'd0 ^ working_key[1322]);
  assign icmp_ln169_fu_860_p2 = ((((working_key[1320] == 1'b1)? rows_1_reg_391 == Const_401 : rows_1_reg_391 > Const_401) ^ working_key[1323]) == 1'b1)? Const_403 : Const_402;
  assign Const_404 = (4'd8 ^ working_key[1327:1324]);
  assign Const_405 = (1'd1 ^ working_key[1329]);
  assign Const_406 = (1'd0 ^ working_key[1330]);
  assign icmp_ln18_fu_1001_p2 = ((((working_key[1328] == 1'b1)? ii_0_i_i_reg_425 == Const_404 : ii_0_i_i_reg_425 != Const_404) ^ working_key[1331]) == 1'b1)? Const_406 : Const_405;
  assign Const_407 = (1'd0 ^ working_key[1333]);
  assign Const_408 = (1'd0 ^ working_key[1334]);
  assign icmp_ln20_fu_1031_p2 = ((((working_key[1332] == 1'b1)? jj_0_i_i_reg_436 === select_ln40_reg_1685 : jj_0_i_i_reg_436 < select_ln40_reg_1685) ^ working_key[1335]) == 1'b1)? Const_408 : Const_407;
  assign Const_409 = (3'd2 ^ working_key[1338:1336]);
  assign Const_410 = (1'd1 ^ working_key[1340]);
  assign Const_411 = (1'd1 ^ working_key[1341]);
  assign icmp_ln34_fu_886_p2 = ((((working_key[1339] == 1'b1)? i_0_i_reg_402 < Const_409 : i_0_i_reg_402 == Const_409) ^ working_key[1342]) == 1'b1)? Const_410 : Const_411;
  assign Const_412 = (2'd1 ^ working_key[1344:1343]);
  assign Const_413 = (1'd0 ^ working_key[1346]);
  assign Const_414 = (1'd1 ^ working_key[1347]);
  assign icmp_ln39_fu_917_p2 = ((((working_key[1345] == 1'b1)? i_1_i_reg_414 == Const_412 : i_1_i_reg_414 != Const_412) ^ working_key[1348]) == 1'b1)? Const_414 : Const_413;
  assign Const_415 = (4'd15 ^ working_key[1352:1349]);
  assign Const_416 = (1'd1 ^ working_key[1354]);
  assign Const_417 = (1'd1 ^ working_key[1355]);
  assign icmp_ln51_fu_1174_p2 = ((((working_key[1353] == 1'b1)? i_0_i_i_reg_481 == Const_415 : i_0_i_i_reg_481 === Const_415) ^ working_key[1356]) == 1'b1)? Const_416 : Const_417;
  assign Const_418 = (4'd0 ^ working_key[1360:1357]);
  assign Const_419 = (1'd0 ^ working_key[1362]);
  assign Const_420 = (1'd0 ^ working_key[1363]);
  assign icmp_ln70_fu_1239_p2 = ((((working_key[1361] == 1'b1)? jj_0_i_i21_0_reg_492 > Const_418 : jj_0_i_i21_0_reg_492 == Const_418) ^ working_key[1364]) == 1'b1)? Const_420 : Const_419;
  assign Const_421 = (4'd0 ^ working_key[1368:1365]);
  assign Const_422 = (1'd0 ^ working_key[1370]);
  assign Const_423 = (1'd0 ^ working_key[1371]);
  assign icmp_ln72_fu_1301_p2 = ((((working_key[1369] == 1'b1)? kk_0_i_i_0_reg_503 > Const_421 : kk_0_i_i_0_reg_503 == Const_421) ^ working_key[1372]) == 1'b1)? Const_423 : Const_422;
  assign Const_424 = (2'd3 ^ working_key[1374:1373]);
  assign Const_425 = (1'd0 ^ working_key[1376]);
  assign Const_426 = (1'd0 ^ working_key[1377]);
  assign icmp_ln87_1_fu_1428_p2 = ((((working_key[1375] == 1'b1)? level_assign_reg_526 === Const_424 : level_assign_reg_526 == Const_424) ^ working_key[1378]) == 1'b1)? Const_425 : Const_426;
  assign Const_427 = (1'd1 ^ working_key[1380]);
  assign Const_428 = (1'd0 ^ working_key[1381]);
  assign icmp_ln87_fu_1442_p2 = ((((working_key[1379] == 1'b1)? ii_0_i_i25_reg_537 != select_ln87_reg_1885 : ii_0_i_i25_reg_537 < select_ln87_reg_1885) ^ working_key[1382]) == 1'b1)? Const_428 : Const_427;
  assign Const_429 = (4'd0 ^ working_key[1386:1383]);
  assign Const_430 = (1'd0 ^ working_key[1388]);
  assign Const_431 = (1'd0 ^ working_key[1389]);
  assign icmp_ln88_fu_1524_p2 = ((((working_key[1387] == 1'b1)? jj_0_i10_i_reg_548 === Const_429 : jj_0_i10_i_reg_548 == Const_429) ^ working_key[1390]) == 1'b1)? Const_431 : Const_430;
  assign Const_432 = (4'd11 ^ working_key[1394:1391]);
  assign ii_1_fu_1447_p2 = (working_key[1395] == 1'b1)? ii_0_i_i25_reg_537 >> Const_432 : ii_0_i_i25_reg_537 + Const_432;
  assign Const_433 = (4'd4 ^ working_key[1399:1396]);
  assign ii_fu_1007_p2 = (working_key[1400] == 1'b1)? ii_0_i_i_reg_425 + Const_433 : ii_0_i_i_reg_425 * Const_433;
  assign inputs_address0 = zext_ln35_2_fu_907_p1;
  assign Const_434 = (2'd1 ^ working_key[1402:1401]);
  assign j_2_fu_1362_p2 = (working_key[1403] == 1'b1)? level_assign_reg_526 * Const_434 : level_assign_reg_526 + Const_434;
  assign Const_435 = (4'd7 ^ working_key[1407:1404]);
  assign j_fu_1154_p2 = (working_key[1408] == 1'b1)? j_0_i_reg_470 * Const_435 : j_0_i_reg_470 + Const_435;
  assign Const_436 = (7'd84 ^ working_key[1415:1409]);
  assign jj_1_fu_770_p2 = (working_key[1416] == 1'b1)? jj_0_reg_368 + Const_436 : jj_0_reg_368 >> Const_436;
  assign Const_437 = (4'd11 ^ working_key[1420:1417]);
  assign jj_2_fu_1530_p2 = (working_key[1421] == 1'b1)? jj_0_i10_i_reg_548 >> Const_437 : jj_0_i10_i_reg_548 + Const_437;
  assign Const_438 = (4'd3 ^ working_key[1425:1422]);
  assign jj_fu_1036_p2 = (working_key[1426] == 1'b1)? jj_0_i_i_reg_436 + Const_438 : jj_0_i_i_reg_436 * Const_438;
  assign p_shl6_cast_fu_1472_p3 = { { add_ln90_2_reg_1898 }, { 3'd0 } };
  assign p_shl_cast_fu_1056_p3 = { { add_ln21_1_fu_1046_p2 }, { 3'd0 } };
  assign Const_439 = (4'd11 ^ working_key[1430:1427]);
  assign rows_2_fu_866_p2 = (working_key[1431] == 1'b1)? rows_1_reg_391 - Const_439 : rows_1_reg_391 + Const_439;
  assign Const_440 = (4'd2 ^ working_key[1435:1432]);
  assign rows_fu_676_p2 = (working_key[1436] == 1'b1)? rows_0_reg_335 + Const_440 : rows_0_reg_335 << Const_440;
  assign Const_441 = (1'd1 ^ working_key[1437]);
  assign Const_442 = (4'd1 ^ working_key[1442:1439]);
  assign Const_443 = (4'd14 ^ working_key[1446:1443]);
  assign select_ln40_fu_963_p3 = ((((working_key[1438] == 1'b1)? trunc_ln40_fu_959_p1[0:0] === Const_441 : trunc_ln40_fu_959_p1[0:0] > Const_441) ^ working_key[1447]) == 1'b1)? Const_442 : Const_443;
  assign Const_444 = (1'd0 ^ working_key[1448]);
  assign Const_445 = (4'd14 ^ working_key[1453:1450]);
  assign Const_446 = (4'd14 ^ working_key[1457:1454]);
  assign select_ln87_fu_1434_p3 = ((((working_key[1449] == 1'b1)? icmp_ln87_1_fu_1428_p2[0:0] === Const_444 : icmp_ln87_1_fu_1428_p2[0:0] != Const_444) ^ working_key[1458]) == 1'b1)? Const_445 : Const_446;
  assign targets_address0 = zext_ln52_5_fu_1199_p1;
  assign tmp_19_fu_652_p3 = { { ee_0_reg_324 }, { 1'd0 } };
  assign tmp_20_fu_696_p3 = { { add_ln160_1_fu_686_p2 }, { 3'd0 } };
  assign tmp_21_fu_708_p3 = { { add_ln160_1_fu_686_p2 }, { 1'd0 } };
  assign tmp_22_fu_818_p3 = { { jj_0_reg_368 }, { 2'd0 } };
  assign tmp_23_fu_830_p3 = { { jj_0_reg_368 }, { 3'd0 } };
  assign tmp_24_fu_842_p3 = { { jj_0_reg_368 }, { 1'd0 } };
  assign tmp_25_fu_788_p3 = { { cols_1_reg_380 }, { 3'd0 } };
  assign tmp_26_fu_800_p3 = { { cols_1_reg_380 }, { 1'd0 } };
  assign tmp_27_fu_929_p3 = { { i_1_i_reg_414 }, { 3'd0 } };
  assign tmp_28_fu_941_p3 = { { i_1_i_reg_414 }, { 1'd0 } };
  assign tmp_29_fu_971_p3 = { { i_1_fu_923_p2 }, { 3'd0 } };
  assign tmp_30_fu_983_p3 = { { i_1_fu_923_p2 }, { 1'd0 } };
  assign tmp_31_fu_1118_p3 = { { i_0_i13_reg_459 }, { 3'd0 } };
  assign tmp_32_fu_1130_p3 = { { i_0_i13_reg_459 }, { 1'd0 } };
  assign tmp_33_fu_1064_p3 = { { add_ln21_1_fu_1046_p2 }, { 1'd0 } };
  assign tmp_34_fu_1271_p3 = { { add_ln73_fu_1260_p2 }, { 3'd0 } };
  assign tmp_35_fu_1283_p3 = { { add_ln73_fu_1260_p2 }, { 1'd0 } };
  assign tmp_36_fu_1368_p3 = { { j_2_fu_1362_p2 }, { 3'd0 } };
  assign tmp_37_fu_1380_p3 = { { j_2_fu_1362_p2 }, { 1'd0 } };
  assign tmp_38_fu_1398_p3 = { { level_assign_reg_526 }, { 3'd0 } };
  assign tmp_39_fu_1410_p3 = { { level_assign_reg_526 }, { 1'd0 } };
  assign tmp_40_fu_1479_p3 = { { add_ln90_2_reg_1898 }, { 1'd0 } };
  assign tmp_41_fu_1496_p3 = { { add_ln90_4_reg_1904 }, { 3'd0 } };
  assign tmp_42_fu_1507_p3 = { { add_ln90_4_reg_1904 }, { 1'd0 } };
  assign tmp_fu_640_p3 = { { ee_0_reg_324 }, { 3'd0 } };
  assign trunc_ln40_fu_959_p1 = i_1_i_reg_414[0:0];
  assign weights_d0 = reg_609;
  assign Const_447 = (64'd3073753658154284245 ^ working_key[1522:1459]);
  assign xor_ln7_1_fu_1096_p2 = (working_key[1523] == 1'b1)? bitcast_ln7_2_fu_1092_p1 & Const_447 : bitcast_ln7_2_fu_1092_p1 ^ Const_447;
  assign Const_448 = (64'd1348086146912679509 ^ working_key[1587:1524]);
  assign xor_ln7_2_fu_1346_p2 = (working_key[1588] == 1'b1)? bitcast_ln7_4_fu_1342_p1 & Const_448 : bitcast_ln7_4_fu_1342_p1 ^ Const_448;
  assign Const_449 = (64'd3074281423752265013 ^ working_key[1652:1589]);
  assign xor_ln7_fu_1219_p2 = (working_key[1653] == 1'b1)? bitcast_ln7_fu_1215_p1 << Const_449 : bitcast_ln7_fu_1215_p1 ^ Const_449;
  assign zext_ln112_1_fu_1138_p1 = tmp_32_fu_1130_p3;
  assign zext_ln112_2_fu_1160_p1 = j_0_i_reg_470;
  assign zext_ln112_3_fu_1169_p1 = add_ln112_1_fu_1164_p2;
  assign zext_ln112_fu_1126_p1 = tmp_31_fu_1118_p3;
  assign zext_ln160_1_fu_660_p1 = tmp_19_fu_652_p3;
  assign zext_ln160_2_fu_682_p1 = rows_0_reg_335;
  assign zext_ln160_3_fu_691_p1 = add_ln160_1_fu_686_p2;
  assign zext_ln160_4_fu_704_p1 = tmp_20_fu_696_p3;
  assign zext_ln160_5_fu_716_p1 = tmp_21_fu_708_p3;
  assign zext_ln160_6_fu_738_p1 = cols_0_reg_346;
  assign zext_ln160_7_fu_747_p1 = add_ln160_3_fu_742_p2;
  assign zext_ln160_fu_648_p1 = tmp_fu_640_p3;
  assign zext_ln170_1_fu_808_p1 = tmp_26_fu_800_p3;
  assign zext_ln170_2_fu_872_p1 = rows_1_reg_391;
  assign zext_ln170_3_fu_881_p1 = add_ln170_1_fu_876_p2;
  assign zext_ln170_fu_796_p1 = tmp_25_fu_788_p3;
  assign zext_ln21_1_fu_949_p1 = tmp_28_fu_941_p3;
  assign zext_ln21_2_fu_1042_p1 = jj_0_i_i_reg_436;
  assign zext_ln21_3_fu_1051_p1 = add_ln21_1_fu_1046_p2;
  assign zext_ln21_4_fu_1072_p1 = tmp_33_fu_1064_p3;
  assign zext_ln21_5_fu_1087_p1 = add_ln21_3_fu_1082_p2;
  assign zext_ln21_fu_937_p1 = tmp_27_fu_929_p3;
  assign zext_ln23_1_fu_991_p1 = tmp_30_fu_983_p3;
  assign zext_ln23_2_fu_1013_p1 = ii_0_i_i_reg_425;
  assign zext_ln23_3_fu_1017_p1 = ii_0_i_i_reg_425;
  assign zext_ln23_4_fu_1026_p1 = add_ln23_1_fu_1021_p2;
  assign zext_ln23_fu_979_p1 = tmp_29_fu_971_p3;
  assign zext_ln35_1_fu_898_p1 = i_0_i_reg_402;
  assign zext_ln35_2_fu_907_p1 = add_ln35_fu_902_p2;
  assign zext_ln35_fu_912_p1 = i_0_i_reg_402;
  assign zext_ln52_1_fu_838_p1 = tmp_23_fu_830_p3;
  assign zext_ln52_2_fu_850_p1 = tmp_24_fu_842_p3;
  assign zext_ln52_3_fu_1186_p1 = i_0_i_i_reg_481;
  assign zext_ln52_4_fu_1190_p1 = i_0_i_i_reg_481;
  assign zext_ln52_5_fu_1199_p1 = add_ln52_1_fu_1194_p2;
  assign zext_ln52_6_fu_1210_p1 = add_ln52_2_fu_1204_p2;
  assign zext_ln52_fu_826_p1 = tmp_22_fu_818_p3;
  assign zext_ln53_fu_1234_p1 = add_ln53_fu_1229_p2;
  assign zext_ln73_1_fu_1256_p1 = jj_0_i_i21_0_reg_492;
  assign zext_ln73_2_fu_1266_p1 = add_ln73_fu_1260_p2;
  assign zext_ln73_3_fu_1279_p1 = tmp_34_fu_1271_p3;
  assign zext_ln73_4_fu_1291_p1 = tmp_35_fu_1283_p3;
  assign zext_ln73_5_fu_1313_p1 = kk_0_i_i_0_reg_503;
  assign zext_ln73_6_fu_1317_p1 = kk_0_i_i_0_reg_503;
  assign zext_ln73_7_fu_1326_p1 = add_ln73_2_fu_1321_p2;
  assign zext_ln73_8_fu_1337_p1 = add_ln73_3_fu_1331_p2;
  assign zext_ln73_fu_1251_p1 = jj_0_i_i21_0_reg_492;
  assign zext_ln89_fu_1563_p1 = add_ln89_fu_1558_p2;
  assign zext_ln90_10_fu_1540_p1 = jj_0_i10_i_reg_548;
  assign zext_ln90_11_fu_1544_p1 = jj_0_i10_i_reg_548;
  assign zext_ln90_12_fu_1553_p1 = add_ln90_6_fu_1548_p2;
  assign zext_ln90_13_fu_1573_p1 = add_ln90_7_fu_1568_p2;
  assign zext_ln90_1_fu_1388_p1 = tmp_37_fu_1380_p3;
  assign zext_ln90_2_fu_1406_p1 = tmp_38_fu_1398_p3;
  assign zext_ln90_3_fu_1418_p1 = tmp_39_fu_1410_p3;
  assign zext_ln90_4_fu_1453_p1 = ii_0_i_i25_reg_537;
  assign zext_ln90_5_fu_1462_p1 = add_ln90_2_fu_1457_p2;
  assign zext_ln90_6_fu_1486_p1 = tmp_40_fu_1479_p3;
  assign zext_ln90_7_fu_1503_p1 = tmp_41_fu_1496_p3;
  assign zext_ln90_8_fu_1514_p1 = tmp_42_fu_1507_p3;
  assign zext_ln90_9_fu_1536_p1 = jj_0_i10_i_reg_548;
  assign zext_ln90_fu_1376_p1 = tmp_36_fu_1368_p3;

  always @(posedge ap_clk) begin
    add_ln160_reg_1586[0] <= 1'b0;
    add_ln160_2_reg_1599[0] <= 1'b0;
    add_ln170_reg_1636[0] <= 1'b0;
    zext_ln52_reg_1641[1:0] <= 2'b00;
    zext_ln52_reg_1641[9] <= 1'b0;
    add_ln52_reg_1646[0] <= 1'b0;
    add_ln21_reg_1680[0] <= 1'b0;
    select_ln40_reg_1685[0] <= 1'b0;
    add_ln23_reg_1690[0] <= 1'b0;
    zext_ln23_2_reg_1703[8:4] <= 5'b00000;
    add_ln112_reg_1754[0] <= 1'b0;
    zext_ln52_3_reg_1775[4] <= 1'b0;
    add_ln73_1_reg_1818[0] <= 1'b0;
    deltas_addr_2_reg_1823[4] <= 1'b0;
    add_ln90_reg_1874[0] <= 1'b0;
    add_ln90_1_reg_1880[0] <= 1'b0;
    select_ln87_reg_1885[0] <= 1'b0;
    add_ln90_3_reg_1915[0] <= 1'b0;
    add_ln90_5_reg_1920[0] <= 1'b0;
  end

  assign working_key = { locking_key[1653:0] };

endmodule

